* NGSPICE file created from CompBlock.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

.subckt CompBlock vdd gnd clk vertices[0] vertices[1] vertices[2] vertices[3] vertices[4]
+ vertices[5] vertices[6] vertices[7] vertices[8] vertices[9] vertices[10] vertices[11]
+ vertices[12] vertices[13] vertices[14] vertices[15] cos_alpha[0] cos_alpha[1] cos_alpha[2]
+ cos_alpha[3] cos_alpha[4] cos_alpha[5] cos_alpha[6] cos_alpha[7] cos_alpha[8] cos_alpha[9]
+ cos_alpha[10] cos_alpha[11] cos_alpha[12] cos_alpha[13] cos_alpha[14] cos_alpha[15]
+ sin_alpha[0] sin_alpha[1] sin_alpha[2] sin_alpha[3] sin_alpha[4] sin_alpha[5] sin_alpha[6]
+ sin_alpha[7] sin_alpha[8] sin_alpha[9] sin_alpha[10] sin_alpha[11] sin_alpha[12]
+ sin_alpha[13] sin_alpha[14] sin_alpha[15] cos_beta[0] cos_beta[1] cos_beta[2] cos_beta[3]
+ cos_beta[4] cos_beta[5] cos_beta[6] cos_beta[7] cos_beta[8] cos_beta[9] cos_beta[10]
+ cos_beta[11] cos_beta[12] cos_beta[13] cos_beta[14] cos_beta[15] sin_beta[0] sin_beta[1]
+ sin_beta[2] sin_beta[3] sin_beta[4] sin_beta[5] sin_beta[6] sin_beta[7] sin_beta[8]
+ sin_beta[9] sin_beta[10] sin_beta[11] sin_beta[12] sin_beta[13] sin_beta[14] sin_beta[15]
+ cos_gamma[0] cos_gamma[1] cos_gamma[2] cos_gamma[3] cos_gamma[4] cos_gamma[5] cos_gamma[6]
+ cos_gamma[7] cos_gamma[8] cos_gamma[9] cos_gamma[10] cos_gamma[11] cos_gamma[12]
+ cos_gamma[13] cos_gamma[14] cos_gamma[15] sin_gamma[0] sin_gamma[1] sin_gamma[2]
+ sin_gamma[3] sin_gamma[4] sin_gamma[5] sin_gamma[6] sin_gamma[7] sin_gamma[8] sin_gamma[9]
+ sin_gamma[10] sin_gamma[11] sin_gamma[12] sin_gamma[13] sin_gamma[14] sin_gamma[15]
+ dx[0] dx[1] dx[2] dx[3] dx[4] dx[5] dx[6] dx[7] dx[8] dx[9] dx[10] dx[11] dx[12]
+ dx[13] dx[14] dx[15] dy[0] dy[1] dy[2] dy[3] dy[4] dy[5] dy[6] dy[7] dy[8] dy[9]
+ dy[10] dy[11] dy[12] dy[13] dy[14] dy[15] dz[0] dz[1] dz[2] dz[3] dz[4] dz[5] dz[6]
+ dz[7] dz[8] dz[9] dz[10] dz[11] dz[12] dz[13] dz[14] dz[15] vertices_out[0] vertices_out[1]
+ vertices_out[2] vertices_out[3] vertices_out[4] vertices_out[5] vertices_out[6]
+ vertices_out[7] vertices_out[8] vertices_out[9] vertices_out[10] vertices_out[11]
+ vertices_out[12] vertices_out[13] vertices_out[14] vertices_out[15]
XFILL_22_0_2 gnd vdd FILL
XFILL_5_1_2 gnd vdd FILL
XOAI21X1_382 OR2X2_48/B OR2X2_48/A OAI21X1_382/C gnd INVX1_311/A vdd OAI21X1
XOAI21X1_360 OAI21X1_361/A OAI21X1_361/B INVX1_271/Y gnd OAI21X1_360/Y vdd OAI21X1
XOAI21X1_371 INVX1_226/Y INVX1_18/Y INVX1_304/Y gnd AND2X2_86/A vdd OAI21X1
XAND2X2_5 AND2X2_5/A AND2X2_7/A gnd AND2X2_5/Y vdd AND2X2
XFILL_13_0_2 gnd vdd FILL
XOAI21X1_393 AND2X2_75/Y INVX1_285/Y INVX1_286/Y gnd INVX1_316/A vdd OAI21X1
XINVX1_232 INVX1_232/A gnd INVX1_232/Y vdd INVX1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_210 vertices[10] gnd OAI22X1_9/D vdd INVX1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XOAI21X1_190 AOI21X1_87/Y AOI21X1_88/Y AOI22X1_24/Y gnd AOI21X1_90/A vdd OAI21X1
XINVX1_276 INVX1_276/A gnd INVX1_276/Y vdd INVX1
XINVX1_287 NOR3X1_27/A gnd INVX1_287/Y vdd INVX1
XINVX1_298 cos_gamma[13] gnd INVX1_298/Y vdd INVX1
XINVX1_265 INVX1_265/A gnd INVX1_265/Y vdd INVX1
XNAND2X1_43 INVX1_49/A NAND2X1_43/B gnd NAND3X1_6/C vdd NAND2X1
XNAND2X1_10 BUFX2_3/Y vertices[2] gnd OR2X2_3/B vdd NAND2X1
XNAND2X1_21 cos_gamma[3] INVX1_9/A gnd NOR2X1_43/A vdd NAND2X1
XNAND2X1_32 cos_gamma[3] INVX1_27/Y gnd OAI21X1_36/A vdd NAND2X1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XNAND2X1_98 INVX1_93/Y NOR2X1_64/Y gnd NAND2X1_99/B vdd NAND2X1
XNAND2X1_76 INVX1_87/Y NAND2X1_76/B gnd AOI22X1_4/A vdd NAND2X1
XNAND2X1_87 AND2X2_22/Y AND2X2_23/Y gnd NAND3X1_47/C vdd NAND2X1
XNAND2X1_65 INVX1_15/A vertices[3] gnd INVX1_74/A vdd NAND2X1
XNAND2X1_54 cos_gamma[4] INVX1_18/A gnd OR2X2_13/B vdd NAND2X1
XAOI21X1_247 NAND3X1_516/C OAI21X1_490/Y INVX1_376/A gnd OAI21X1_495/B vdd AOI21X1
XAOI21X1_236 OAI21X1_466/Y NAND3X1_497/A NAND3X1_498/A gnd OAI21X1_511/A vdd AOI21X1
XAOI21X1_258 INVX1_363/A NAND3X1_492/B OAI21X1_467/A gnd NOR3X1_48/B vdd AOI21X1
XAOI21X1_225 NAND3X1_475/Y NAND3X1_476/Y INVX1_357/A gnd OAI21X1_457/B vdd AOI21X1
XAOI21X1_214 OAI21X1_415/Y NAND3X1_450/B INVX1_329/A gnd NOR3X1_43/C vdd AOI21X1
XAOI21X1_203 OAI21X1_398/Y NAND3X1_414/B INVX1_321/Y gnd NOR3X1_38/B vdd AOI21X1
XAOI22X1_41 AOI22X1_41/A AOI22X1_41/B AND2X2_78/Y AOI22X1_41/D gnd AOI22X1_41/Y vdd
+ AOI22X1
XAOI22X1_30 AOI22X1_30/A OR2X2_17/Y AOI22X1_30/C AOI22X1_30/D gnd AOI22X1_30/Y vdd
+ AOI22X1
XAOI22X1_52 INVX1_263/A INVX1_262/Y AND2X2_96/B AOI22X1_52/D gnd NOR3X1_43/B vdd AOI22X1
XNAND3X1_229 OAI21X1_230/Y NAND3X1_232/A INVX1_211/Y gnd OAI21X1_276/C vdd NAND3X1
XNAND3X1_218 NOR2X1_84/Y AND2X2_57/B OAI21X1_203/Y gnd INVX1_192/A vdd NAND3X1
XNAND3X1_207 INVX1_184/Y AND2X2_48/B AOI21X1_99/B gnd AND2X2_48/A vdd NAND3X1
XOAI22X1_3 INVX1_8/Y INVX1_43/Y INVX1_7/Y OAI22X1_8/B gnd OAI22X1_3/Y vdd OAI22X1
XNAND2X1_409 NAND3X1_423/Y NAND3X1_426/Y gnd INVX1_323/A vdd NAND2X1
XFILL_20_1_0 gnd vdd FILL
XAND2X2_110 OR2X2_55/Y AOI22X1_59/B gnd NOR3X1_51/A vdd AND2X2
XFILL_28_2_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 INVX1_19/Y NOR2X1_20/A INVX1_20/A gnd XNOR2X1_8/B vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XNAND2X1_228 XOR2X1_13/Y INVX1_206/Y gnd NAND3X1_234/C vdd NAND2X1
XNAND2X1_217 NAND2X1_217/A NAND3X1_210/B gnd INVX1_221/A vdd NAND2X1
XNAND2X1_206 AND2X2_59/A OR2X2_25/Y gnd NAND3X1_267/A vdd NAND2X1
XNAND2X1_239 AOI22X1_32/A AOI22X1_32/B gnd OAI21X1_242/C vdd NAND2X1
XOR2X2_55 OR2X2_55/A OR2X2_55/B gnd OR2X2_55/Y vdd OR2X2
XOR2X2_33 OR2X2_33/A OR2X2_33/B gnd OR2X2_33/Y vdd OR2X2
XNAND3X1_390 INVX1_258/Y AND2X2_95/B OAI21X1_364/Y gnd AND2X2_95/A vdd NAND3X1
XOR2X2_44 OR2X2_44/A OR2X2_44/B gnd OR2X2_44/Y vdd OR2X2
XOR2X2_11 OR2X2_11/A OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_22 OR2X2_22/A OR2X2_22/B gnd OR2X2_22/Y vdd OR2X2
XXNOR2X1_6 XNOR2X1_6/A XNOR2X1_6/B gnd OR2X2_5/A vdd XNOR2X1
XFILL_25_0_0 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_8_1_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_383 INVX1_29/Y INVX1_203/Y OAI21X1_486/A gnd OAI21X1_384/C vdd OAI21X1
XOAI21X1_350 OAI21X1_379/B NOR3X1_35/Y INVX1_276/A gnd OAI21X1_350/Y vdd OAI21X1
XOAI21X1_361 OAI21X1_361/A OAI21X1_361/B INVX1_271/A gnd AOI22X1_42/D vdd OAI21X1
XOAI21X1_394 INVX1_73/Y NOR2X1_86/B OR2X2_39/A gnd OAI21X1_394/Y vdd OAI21X1
XOAI21X1_372 NOR2X1_133/A NOR2X1_166/A AND2X2_70/B gnd XNOR2X1_41/B vdd OAI21X1
XAND2X2_6 INVX1_24/Y AND2X2_6/B gnd XOR2X1_4/B vdd AND2X2
XXOR2X1_50 XOR2X1_50/A XOR2X1_50/B gnd XOR2X1_50/Y vdd XOR2X1
XINVX1_277 cos_alpha[12] gnd INVX1_277/Y vdd INVX1
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XINVX1_266 INVX1_266/A gnd INVX1_266/Y vdd INVX1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XAOI22X1_1 INVX1_42/A OAI22X1_3/Y INVX1_67/Y INVX1_68/Y gnd OR2X2_8/A vdd AOI22X1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XOAI21X1_191 AOI21X1_91/Y AOI21X1_90/Y AOI21X1_89/Y gnd AOI21X1_92/A vdd OAI21X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XOAI21X1_180 INVX1_45/Y NOR2X1_86/B OR2X2_22/A gnd OAI21X1_180/Y vdd OAI21X1
XINVX1_288 NOR3X1_27/B gnd INVX1_288/Y vdd INVX1
XINVX1_299 INVX1_299/A gnd INVX1_299/Y vdd INVX1
XNAND2X1_44 NAND3X1_8/B NAND3X1_8/A gnd NAND2X1_45/B vdd NAND2X1
XNAND2X1_33 NOR2X1_34/A NOR2X1_34/B gnd NAND2X1_34/A vdd NAND2X1
XNAND2X1_55 OAI21X1_37/Y OAI21X1_62/C gnd OR2X2_8/B vdd NAND2X1
XNAND2X1_22 cos_gamma[2] INVX1_27/Y gnd XNOR2X1_6/B vdd NAND2X1
XNAND2X1_66 BUFX2_2/Y vertices[4] gnd INVX1_102/A vdd NAND2X1
XNAND2X1_11 BUFX2_16/Y vertices[2] gnd OAI21X1_7/B vdd NAND2X1
XNAND2X1_77 cos_gamma[6] INVX1_9/A gnd NOR2X1_82/A vdd NAND2X1
XFILL_28_1 gnd vdd FILL
XNAND2X1_99 OAI21X1_84/Y NAND2X1_99/B gnd OR2X2_12/A vdd NAND2X1
XNAND2X1_88 BUFX2_11/Y vertices[4] gnd INVX1_100/A vdd NAND2X1
XAOI21X1_259 NAND3X1_538/C INVX1_380/Y INVX1_381/Y gnd OAI21X1_509/A vdd AOI21X1
XAOI22X1_53 AOI22X1_53/A AOI22X1_53/B AOI22X1_53/C AOI22X1_53/D gnd NOR3X1_44/B vdd
+ AOI22X1
XAOI21X1_237 NAND3X1_497/Y NAND3X1_498/Y OAI21X1_511/B gnd OAI21X1_471/A vdd AOI21X1
XAOI21X1_248 NAND3X1_468/C NAND3X1_468/B INVX1_354/A gnd OAI21X1_497/A vdd AOI21X1
XAOI21X1_215 AOI21X1_215/A OAI21X1_417/Y NOR3X1_43/Y gnd AOI22X1_56/D vdd AOI21X1
XAOI21X1_226 NAND3X1_426/B NAND3X1_426/C NAND3X1_423/A gnd AOI21X1_227/C vdd AOI21X1
XAOI21X1_204 AND2X2_74/Y OAI21X1_344/Y NOR3X1_31/C gnd NOR3X1_39/A vdd AOI21X1
XAOI22X1_42 AND2X2_84/A AND2X2_81/B AND2X2_93/B AOI22X1_42/D gnd AOI22X1_42/Y vdd
+ AOI22X1
XAOI22X1_20 AOI22X1_20/A AOI22X1_20/B AOI22X1_20/C AOI22X1_20/D gnd AOI22X1_20/Y vdd
+ AOI22X1
XAOI22X1_31 AOI22X1_31/A AOI22X1_31/B INVX1_217/Y AOI22X1_31/D gnd INVX1_237/A vdd
+ AOI22X1
XNAND3X1_219 INVX1_191/A INVX1_192/A OAI21X1_204/Y gnd NAND3X1_275/A vdd NAND3X1
XNAND3X1_208 XOR2X1_11/Y AND2X2_48/A NAND3X1_208/C gnd NAND3X1_210/B vdd NAND3X1
XOAI22X1_4 INVX1_16/Y INVX1_46/Y INVX1_29/Y INVX1_28/Y gnd OAI22X1_4/Y vdd OAI22X1
XFILL_20_1_1 gnd vdd FILL
XAND2X2_100 AND2X2_100/A AND2X2_100/B gnd AND2X2_100/Y vdd AND2X2
XFILL_28_2_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XNAND2X1_229 NAND3X1_226/Y NAND3X1_227/Y gnd NAND3X1_237/C vdd NAND2X1
XNAND2X1_207 AND2X2_53/B AND2X2_53/A gnd OAI21X1_247/C vdd NAND2X1
XNAND2X1_218 cos_gamma[2] NAND3X1_457/B gnd INVX1_217/A vdd NAND2X1
XNAND3X1_391 NAND3X1_391/A AND2X2_94/A INVX1_296/Y gnd NAND3X1_395/B vdd NAND3X1
XNAND3X1_380 NAND3X1_380/A AND2X2_92/B NAND3X1_380/C gnd AND2X2_92/A vdd NAND3X1
XFILL_10_1 gnd vdd FILL
XOR2X2_34 OR2X2_34/A OR2X2_34/B gnd OR2X2_34/Y vdd OR2X2
XOR2X2_45 OR2X2_45/A OR2X2_45/B gnd OR2X2_45/Y vdd OR2X2
XOR2X2_56 OR2X2_56/A OR2X2_56/B gnd OR2X2_56/Y vdd OR2X2
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 XNOR2X1_7/A INVX1_32/Y gnd XNOR2X1_8/A vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XOAI21X1_510 NOR3X1_48/A NOR3X1_48/C NOR3X1_48/B gnd OAI21X1_510/Y vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XOAI21X1_384 XOR2X1_23/B OAI21X1_437/C OAI21X1_384/C gnd OR2X2_38/A vdd OAI21X1
XOAI21X1_395 NOR3X1_27/A NOR3X1_27/B OAI21X1_395/C gnd OAI21X1_395/Y vdd OAI21X1
XOAI21X1_362 AOI22X1_42/Y OAI21X1_363/B OAI21X1_362/C gnd AOI22X1_43/D vdd OAI21X1
XOAI21X1_351 OAI21X1_351/A NOR3X1_34/Y INVX1_291/A gnd AND2X2_79/A vdd OAI21X1
XOAI21X1_340 INVX1_244/A NOR2X1_126/Y OAI21X1_340/C gnd OAI21X1_340/Y vdd OAI21X1
XOAI21X1_373 NOR2X1_83/A INVX1_124/Y NOR2X1_169/A gnd OAI21X1_374/C vdd OAI21X1
XAND2X2_7 AND2X2_7/A OR2X2_3/Y gnd AND2X2_8/B vdd AND2X2
XNAND2X1_390 OAI21X1_385/Y OR2X2_38/Y gnd OAI21X1_432/B vdd NAND2X1
XXOR2X1_40 XOR2X1_40/A XOR2X1_40/B gnd XOR2X1_40/Y vdd XOR2X1
XXOR2X1_51 XOR2X1_51/A XOR2X1_51/B gnd OR2X2_59/A vdd XOR2X1
XAOI22X1_2 INVX1_52/Y AOI22X1_2/B INVX1_51/Y NAND3X1_4/B gnd NOR3X1_1/A vdd AOI22X1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XINVX1_267 INVX1_267/A gnd INVX1_267/Y vdd INVX1
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XINVX1_245 vertices[11] gnd OAI22X1_9/B vdd INVX1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XOAI21X1_170 OR2X2_16/B OR2X2_16/A OR2X2_18/Y gnd INVX1_172/A vdd OAI21X1
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XOAI21X1_192 AOI21X1_91/Y AOI21X1_90/Y OAI21X1_192/C gnd AOI21X1_93/A vdd OAI21X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XINVX1_256 INVX1_256/A gnd INVX1_256/Y vdd INVX1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XOAI21X1_181 NOR2X1_96/Y AND2X2_42/Y INVX1_176/A gnd OAI21X1_181/Y vdd OAI21X1
XNAND2X1_67 OAI21X1_48/Y NAND3X1_18/Y gnd NAND3X1_20/B vdd NAND2X1
XNAND2X1_78 OAI21X1_60/Y INVX1_92/Y gnd INVX1_93/A vdd NAND2X1
XNAND2X1_45 AOI21X1_5/Y NAND2X1_45/B gnd NOR2X1_60/A vdd NAND2X1
XNAND2X1_34 NAND2X1_34/A INVX1_38/Y gnd INVX1_39/A vdd NAND2X1
XNAND2X1_23 cos_gamma[1] INVX1_18/A gnd XNOR2X1_5/B vdd NAND2X1
XNAND2X1_56 OR2X2_8/B OR2X2_8/A gnd NAND3X1_14/B vdd NAND2X1
XNAND2X1_12 NOR2X1_17/A AND2X2_5/Y gnd INVX1_17/A vdd NAND2X1
XNAND2X1_89 BUFX2_17/Y vertices[5] gnd NOR2X1_58/A vdd NAND2X1
XFILL_28_2 gnd vdd FILL
XAOI21X1_205 OAI21X1_400/Y OAI21X1_441/C AND2X2_91/Y gnd NOR3X1_39/B vdd AOI21X1
XAOI21X1_216 INVX1_307/A NAND3X1_436/C NOR2X1_170/Y gnd OR2X2_47/A vdd AOI21X1
XAOI21X1_238 NAND3X1_494/B AOI22X1_60/A XNOR2X1_46/Y gnd OAI21X1_471/B vdd AOI21X1
XAOI21X1_249 INVX1_356/Y OAI21X1_452/Y NOR3X1_44/Y gnd NAND3X1_523/A vdd AOI21X1
XAOI22X1_54 AOI22X1_55/A AOI22X1_55/B AOI22X1_54/C AOI22X1_54/D gnd AOI22X1_54/Y vdd
+ AOI22X1
XAOI21X1_227 INVX1_323/A INVX1_359/Y AOI21X1_227/C gnd OAI21X1_458/C vdd AOI21X1
XAOI22X1_43 INVX1_329/A AOI22X1_43/B AND2X2_94/B AOI22X1_43/D gnd AOI22X1_43/Y vdd
+ AOI22X1
XAOI22X1_21 cos_gamma[2] NOR2X1_73/Y AOI22X1_21/C AOI22X1_21/D gnd NOR3X1_15/B vdd
+ AOI22X1
XAOI22X1_32 AOI22X1_32/A AOI22X1_32/B AOI22X1_32/C AOI22X1_32/D gnd AOI22X1_32/Y vdd
+ AOI22X1
XAOI22X1_10 vertices[0] cos_alpha[7] vertices[1] cos_alpha[6] gnd NOR2X1_75/A vdd
+ AOI22X1
XNAND3X1_209 INVX1_188/A NAND3X1_210/B OAI21X1_198/Y gnd AND2X2_53/B vdd NAND3X1
XOAI22X1_5 OAI22X1_5/A OAI22X1_5/B XOR2X1_9/B XOR2X1_9/A gnd OAI22X1_5/Y vdd OAI22X1
XFILL_20_1_2 gnd vdd FILL
XAND2X2_101 AOI22X1_53/B AOI22X1_53/A gnd AND2X2_101/Y vdd AND2X2
XFILL_28_2_2 gnd vdd FILL
XFILL_3_2_2 gnd vdd FILL
XFILL_11_1_2 gnd vdd FILL
XFILL_19_2_2 gnd vdd FILL
XNAND3X1_540 AOI22X1_59/C INVX1_382/Y AOI22X1_59/D gnd NAND3X1_541/B vdd NAND3X1
XNAND2X1_219 vertices[1] cos_alpha[9] gnd NOR2X1_140/A vdd NAND2X1
XNAND2X1_208 cos_gamma[3] NAND2X1_536/B gnd OAI21X1_263/A vdd NAND2X1
XNAND3X1_392 OR2X2_27/Y NAND3X1_395/B OAI21X1_365/Y gnd NAND3X1_393/C vdd NAND3X1
XNAND3X1_381 INVX1_271/A NAND3X1_383/A AND2X2_92/A gnd NAND3X1_382/A vdd NAND3X1
XNAND3X1_370 INVX1_273/A AND2X2_89/B OAI21X1_356/Y gnd AND2X2_89/A vdd NAND3X1
XOR2X2_35 OR2X2_41/A OR2X2_35/B gnd OR2X2_35/Y vdd OR2X2
XOR2X2_57 OR2X2_57/A OR2X2_57/B gnd OR2X2_57/Y vdd OR2X2
XOR2X2_46 OR2X2_46/A OR2X2_46/B gnd OR2X2_46/Y vdd OR2X2
XOR2X2_24 OR2X2_24/A OR2X2_24/B gnd OR2X2_24/Y vdd OR2X2
XXNOR2X1_8 XNOR2X1_8/A XNOR2X1_8/B gnd OR2X2_5/B vdd XNOR2X1
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XFILL_25_0_2 gnd vdd FILL
XFILL_0_0_2 gnd vdd FILL
XOAI21X1_511 OAI21X1_511/A OAI21X1_511/B AOI22X1_60/A gnd OAI21X1_511/Y vdd OAI21X1
XINVX1_8 cos_gamma[1] gnd INVX1_8/Y vdd INVX1
XOAI21X1_500 INVX1_65/Y NOR2X1_197/B OAI21X1_500/C gnd OAI21X1_500/Y vdd OAI21X1
XFILL_8_1_2 gnd vdd FILL
XFILL_16_0_2 gnd vdd FILL
XFILL_9_1 gnd vdd FILL
XOAI21X1_330 INVX1_279/A INVX1_280/Y OAI21X1_330/C gnd OAI21X1_330/Y vdd OAI21X1
XOAI21X1_341 NOR3X1_27/B NOR3X1_27/C NOR3X1_27/A gnd OAI21X1_341/Y vdd OAI21X1
XOAI21X1_385 INVX1_16/Y INVX1_241/Y OR2X2_38/A gnd OAI21X1_385/Y vdd OAI21X1
XOAI21X1_363 AOI22X1_42/Y OAI21X1_363/B OAI21X1_363/C gnd OAI21X1_363/Y vdd OAI21X1
XOAI21X1_352 NOR3X1_34/B NOR3X1_34/C NOR3X1_34/A gnd OAI21X1_352/Y vdd OAI21X1
XOAI21X1_396 AND2X2_90/Y NOR2X1_160/Y INVX1_318/Y gnd OAI21X1_396/Y vdd OAI21X1
XOAI21X1_374 NOR2X1_166/A NOR2X1_166/B OAI21X1_374/C gnd XNOR2X1_40/A vdd OAI21X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XNAND2X1_391 INVX1_312/A OAI21X1_432/B gnd NAND3X1_402/C vdd NAND2X1
XXOR2X1_52 XOR2X1_52/A XOR2X1_52/B gnd XOR2X1_52/Y vdd XOR2X1
XXOR2X1_30 XOR2X1_30/A XOR2X1_30/B gnd XOR2X1_30/Y vdd XOR2X1
XNAND2X1_380 XOR2X1_24/B XOR2X1_24/A gnd NAND2X1_381/A vdd NAND2X1
XXOR2X1_41 XOR2X1_41/A XOR2X1_41/B gnd XOR2X1_41/Y vdd XOR2X1
XOAI21X1_160 AOI22X1_22/Y AOI21X1_76/Y INVX1_163/Y gnd AOI21X1_77/A vdd OAI21X1
XAOI22X1_3 BUFX2_13/Y vertices[3] AOI22X1_7/D AOI22X1_3/D gnd NOR3X1_1/B vdd AOI22X1
XOAI21X1_171 INVX1_36/Y OAI22X1_8/D OR2X2_19/A gnd OAI21X1_171/Y vdd OAI21X1
XOAI21X1_182 NOR2X1_96/Y AND2X2_42/Y INVX1_176/Y gnd OAI21X1_182/Y vdd OAI21X1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XINVX1_235 INVX1_235/A gnd OR2X2_28/B vdd INVX1
XOAI21X1_193 AOI21X1_92/Y AOI21X1_93/Y OAI21X1_193/C gnd AOI21X1_97/B vdd OAI21X1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XINVX1_213 INVX1_213/A gnd INVX1_213/Y vdd INVX1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XNAND2X1_68 NAND3X1_22/Y NAND3X1_24/Y gnd INVX1_78/A vdd NAND2X1
XNAND2X1_46 NOR2X1_60/A NAND3X1_8/Y gnd OAI22X1_8/B vdd NAND2X1
XNAND2X1_35 XNOR2X1_8/B XNOR2X1_8/A gnd OAI21X1_22/C vdd NAND2X1
XNAND2X1_13 NAND3X1_2/Y OAI21X1_9/Y gnd XOR2X1_1/A vdd NAND2X1
XNAND2X1_57 NAND3X1_14/B OR2X2_8/Y gnd OAI21X1_38/C vdd NAND2X1
XNAND2X1_24 vertices[1] BUFX2_11/Y gnd INVX1_48/A vdd NAND2X1
XNAND2X1_79 cos_gamma[3] INVX1_43/A gnd OR2X2_13/A vdd NAND2X1
XAOI21X1_239 NAND3X1_453/B AND2X2_96/A NAND3X1_453/A gnd OAI21X1_472/A vdd AOI21X1
XAOI21X1_206 OAI21X1_399/Y NAND3X1_416/B OAI21X1_389/Y gnd NOR3X1_40/B vdd AOI21X1
XAOI21X1_217 NAND3X1_440/C AOI22X1_46/D INVX1_340/Y gnd INVX1_341/A vdd AOI21X1
XAOI21X1_228 NAND2X1_411/B NAND3X1_427/Y INVX1_8/Y gnd NAND3X1_484/B vdd AOI21X1
XAOI22X1_44 AOI22X1_44/A AOI22X1_44/B AOI22X1_44/C AOI22X1_44/D gnd NOR2X1_153/A vdd
+ AOI22X1
XAOI22X1_55 AOI22X1_55/A AOI22X1_55/B AOI22X1_55/C AOI22X1_55/D gnd AOI22X1_55/Y vdd
+ AOI22X1
XAOI22X1_33 AND2X2_72/A AOI22X1_33/B INVX1_270/A AOI22X1_33/D gnd AOI22X1_33/Y vdd
+ AOI22X1
XAOI22X1_22 AND2X2_39/A AND2X2_39/B AOI22X1_22/C AOI22X1_22/D gnd AOI22X1_22/Y vdd
+ AOI22X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XAOI22X1_11 INVX1_15/A vertices[5] NAND3X1_71/B NAND3X1_71/C gnd NOR3X1_13/B vdd AOI22X1
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 INVX1_1/Y OAI22X1_6/B INVX1_10/Y OAI22X1_6/D gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XAND2X2_102 AND2X2_102/A AOI22X1_48/C gnd AND2X2_102/Y vdd AND2X2
XNAND3X1_541 NOR2X1_200/A NAND3X1_541/B OAI21X1_512/Y gnd NAND3X1_542/A vdd NAND3X1
XNAND3X1_530 NAND3X1_530/A OAI21X1_501/Y INVX1_378/Y gnd NAND3X1_531/B vdd NAND3X1
XNAND2X1_209 cos_gamma[4] NAND2X1_536/B gnd OR2X2_31/B vdd NAND2X1
XFILL_28_0_0 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_19_0_0 gnd vdd FILL
XNAND3X1_360 OAI21X1_380/C OAI21X1_346/Y INVX1_282/Y gnd NAND3X1_362/C vdd NAND3X1
XNAND3X1_382 NAND3X1_382/A NAND3X1_382/B OAI21X1_360/Y gnd NAND3X1_387/A vdd NAND3X1
XNAND3X1_371 XOR2X1_24/Y AND2X2_89/A NAND3X1_373/C gnd NAND3X1_377/A vdd NAND3X1
XNAND3X1_393 INVX1_297/A AND2X2_95/A NAND3X1_393/C gnd AOI22X1_44/A vdd NAND3X1
XOR2X2_14 OR2X2_14/A OR2X2_14/B gnd OR2X2_14/Y vdd OR2X2
XOR2X2_58 OR2X2_58/A OR2X2_58/B gnd OR2X2_58/Y vdd OR2X2
XOR2X2_47 OR2X2_47/A OR2X2_47/B gnd OR2X2_47/Y vdd OR2X2
XOR2X2_36 OR2X2_36/A OR2X2_36/B gnd OR2X2_36/Y vdd OR2X2
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XXNOR2X1_9 XOR2X1_4/Y XNOR2X1_9/B gnd XNOR2X1_9/Y vdd XNOR2X1
XOR2X2_25 OR2X2_25/A OR2X2_25/B gnd OR2X2_25/Y vdd OR2X2
XOAI21X1_512 NOR3X1_50/A NOR3X1_50/C NOR3X1_50/B gnd OAI21X1_512/Y vdd OAI21X1
XOAI21X1_501 INVX1_22/Y NOR2X1_196/B NOR2X1_198/B gnd OAI21X1_501/Y vdd OAI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND2X1_540 AND2X2_109/B AND2X2_109/A gnd NOR3X1_47/A vdd NAND2X1
XFILL_9_2 gnd vdd FILL
XNAND3X1_190 NAND3X1_190/A OAI21X1_193/C NAND3X1_190/C gnd AOI21X1_96/B vdd NAND3X1
XOAI21X1_342 NOR3X1_29/A NOR3X1_29/C NOR3X1_29/B gnd OAI21X1_342/Y vdd OAI21X1
XOAI21X1_364 AOI22X1_43/Y OAI21X1_365/B INVX1_296/Y gnd OAI21X1_364/Y vdd OAI21X1
XOAI21X1_331 OAI21X1_331/A OAI21X1_331/B OAI21X1_331/C gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_353 OAI21X1_353/A AOI22X1_32/Y AND2X2_64/A gnd OAI21X1_458/A vdd OAI21X1
XOAI21X1_320 OR2X2_28/B OR2X2_28/A OR2X2_31/Y gnd INVX1_272/A vdd OAI21X1
XOAI21X1_386 NOR2X1_143/Y OAI21X1_386/B OAI21X1_386/C gnd INVX1_313/A vdd OAI21X1
XOAI21X1_375 XNOR2X1_38/Y OAI21X1_375/B AND2X2_87/A gnd XNOR2X1_42/A vdd OAI21X1
XXOR2X1_20 XOR2X1_20/A XOR2X1_20/B gnd XOR2X1_20/Y vdd XOR2X1
XOAI21X1_397 INVX1_1/Y INVX1_319/Y OR2X2_40/A gnd OAI21X1_397/Y vdd OAI21X1
XAND2X2_9 AND2X2_9/A INVX1_30/Y gnd AND2X2_9/Y vdd AND2X2
XNAND2X1_392 INVX1_312/Y OAI21X1_432/B gnd NAND3X1_403/C vdd NAND2X1
XXOR2X1_31 XOR2X1_31/A XOR2X1_31/B gnd XOR2X1_31/Y vdd XOR2X1
XXOR2X1_42 dy[15] dz[15] gnd XOR2X1_42/Y vdd XOR2X1
XNAND2X1_370 OAI21X1_418/C NAND2X1_370/B gnd OAI21X1_418/B vdd NAND2X1
XNAND2X1_381 NAND2X1_381/A NAND3X1_377/A gnd INVX1_327/A vdd NAND2X1
XINVX1_203 cos_alpha[10] gnd INVX1_203/Y vdd INVX1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XAOI22X1_4 AOI22X1_4/A NOR3X1_12/A INVX1_61/Y NOR2X1_42/Y gnd NOR2X1_52/A vdd AOI22X1
XOAI21X1_161 NOR3X1_16/B NOR3X1_16/C NOR3X1_16/A gnd AOI21X1_78/A vdd OAI21X1
XOAI21X1_150 AOI22X1_18/Y AOI21X1_66/Y AOI21X1_85/C gnd AOI22X1_20/C vdd OAI21X1
XOAI21X1_194 AOI21X1_92/Y AOI21X1_93/Y AOI21X1_94/Y gnd AOI21X1_96/A vdd OAI21X1
XOAI21X1_172 INVX1_65/Y OAI22X1_8/B OAI21X1_172/C gnd AND2X2_40/A vdd OAI21X1
XOAI21X1_183 AOI21X1_86/Y AOI21X1_66/C INVX1_181/A gnd OAI21X1_192/C vdd OAI21X1
XNAND2X1_14 dy[2] dx[2] gnd INVX1_20/A vdd NAND2X1
XINVX1_258 OR2X2_27/Y gnd INVX1_258/Y vdd INVX1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XNAND2X1_25 BUFX2_17/Y vertices[3] gnd AND2X2_18/A vdd NAND2X1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XNAND2X1_69 INVX1_78/A NOR2X1_48/Y gnd NAND2X1_70/B vdd NAND2X1
XNAND2X1_47 cos_gamma[1] AND2X2_13/Y gnd INVX1_68/A vdd NAND2X1
XNAND2X1_58 AND2X2_19/A OAI21X1_38/Y gnd INVX1_69/A vdd NAND2X1
XNAND2X1_36 AND2X2_8/B AND2X2_8/A gnd AOI21X1_2/B vdd NAND2X1
XAOI21X1_229 NAND3X1_485/B NAND3X1_485/C INVX1_348/A gnd OAI21X1_461/A vdd AOI21X1
XAOI21X1_207 INVX1_282/Y OAI21X1_346/Y NOR3X1_33/C gnd NOR3X1_41/A vdd AOI21X1
XAOI21X1_218 NAND3X1_308/Y OAI21X1_296/Y INVX1_36/Y gnd OAI21X1_500/C vdd AOI21X1
XAOI22X1_12 NAND3X1_70/Y OAI21X1_99/Y NAND3X1_78/A NAND3X1_78/C gnd NOR3X1_14/A vdd
+ AOI22X1
XAOI22X1_23 INVX1_152/Y NOR2X1_77/B NOR2X1_87/Y AOI22X1_23/D gnd INVX1_176/A vdd AOI22X1
XAOI22X1_56 AOI22X1_56/A AOI22X1_56/B AOI22X1_56/C AOI22X1_56/D gnd NOR2X1_179/A vdd
+ AOI22X1
XAOI22X1_45 cos_gamma[2] AOI22X1_45/B AOI22X1_45/C AOI22X1_45/D gnd NOR3X1_42/B vdd
+ AOI22X1
XAOI22X1_34 AOI22X1_34/A AOI22X1_34/B AOI22X1_34/C AOI22X1_34/D gnd AOI22X1_34/Y vdd
+ AOI22X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_7/A OAI22X1_7/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XAND2X2_103 AND2X2_103/A AOI22X1_50/C gnd AND2X2_103/Y vdd AND2X2
XNAND3X1_520 NAND3X1_522/A OAI21X1_495/Y XNOR2X1_77/Y gnd NAND3X1_521/C vdd NAND3X1
XNAND3X1_542 NAND3X1_542/A OAI21X1_513/Y XNOR2X1_83/Y gnd NAND3X1_543/B vdd NAND3X1
XNAND3X1_531 NAND3X1_531/A NAND3X1_531/B OAI21X1_504/Y gnd NAND3X1_532/B vdd NAND3X1
XFILL_28_0_1 gnd vdd FILL
XFILL_3_0_1 gnd vdd FILL
XFILL_19_0_1 gnd vdd FILL
XNAND3X1_350 INVX1_242/A OAI21X1_330/Y NAND3X1_350/C gnd NAND3X1_350/Y vdd NAND3X1
XOR2X2_48 OR2X2_48/A OR2X2_48/B gnd OR2X2_48/Y vdd OR2X2
XNAND3X1_361 OAI21X1_347/Y NAND3X1_362/C OAI21X1_349/C gnd OAI21X1_379/C vdd NAND3X1
XNAND3X1_383 NAND3X1_383/A AND2X2_92/A INVX1_271/Y gnd AND2X2_93/B vdd NAND3X1
XNAND3X1_394 OR2X2_27/Y AND2X2_95/B OAI21X1_364/Y gnd NAND3X1_396/B vdd NAND3X1
XNAND3X1_372 NAND3X1_378/A NAND3X1_377/A OAI21X1_358/Y gnd AND2X2_92/B vdd NAND3X1
XOR2X2_37 OR2X2_37/A OR2X2_37/B gnd OR2X2_37/Y vdd OR2X2
XOR2X2_26 OR2X2_26/A OR2X2_26/B gnd OR2X2_26/Y vdd OR2X2
XOR2X2_15 OR2X2_15/A OR2X2_15/B gnd OR2X2_15/Y vdd OR2X2
XOR2X2_59 OR2X2_59/A OR2X2_59/B gnd OR2X2_59/Y vdd OR2X2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XOAI21X1_513 NOR3X1_51/B NOR3X1_51/C NOR3X1_51/A gnd OAI21X1_513/Y vdd OAI21X1
XOAI21X1_502 OAI21X1_504/A NOR2X1_198/Y INVX1_378/Y gnd OAI21X1_502/Y vdd OAI21X1
XNAND2X1_541 AOI22X1_59/B OR2X2_55/Y gnd NOR2X1_200/A vdd NAND2X1
XNAND2X1_530 OAI21X1_297/Y NAND3X1_311/C gnd OAI21X1_499/B vdd NAND2X1
XNAND3X1_191 AND2X2_45/Y AOI21X1_96/B AOI21X1_96/A gnd NAND3X1_194/B vdd NAND3X1
XNAND3X1_180 NAND3X1_180/A NAND3X1_180/B OAI21X1_189/C gnd INVX1_212/A vdd NAND3X1
XOAI21X1_387 OAI21X1_388/A OAI21X1_388/B INVX1_313/Y gnd OAI21X1_387/Y vdd OAI21X1
XOAI21X1_398 NOR3X1_36/A NOR3X1_36/C XOR2X1_30/Y gnd OAI21X1_398/Y vdd OAI21X1
XOAI21X1_365 AOI22X1_43/Y OAI21X1_365/B INVX1_296/A gnd OAI21X1_365/Y vdd OAI21X1
XOAI21X1_343 NOR3X1_28/B NOR3X1_28/C NOR3X1_28/A gnd OAI21X1_343/Y vdd OAI21X1
XOAI21X1_332 INVX1_177/Y INVX1_148/Y OR2X2_32/A gnd OAI21X1_333/C vdd OAI21X1
XOAI21X1_376 XOR2X1_22/B XOR2X1_22/A OR2X2_37/Y gnd INVX1_307/A vdd OAI21X1
XOAI21X1_321 OR2X2_31/A OAI21X1_377/C OAI21X1_321/C gnd XOR2X1_22/A vdd OAI21X1
XOAI21X1_310 INVX1_225/A OAI21X1_310/B AOI22X1_37/C gnd INVX1_296/A vdd OAI21X1
XOAI21X1_354 OAI21X1_354/A OAI21X1_354/B AND2X2_78/Y gnd OAI21X1_354/Y vdd OAI21X1
XXOR2X1_32 XOR2X1_32/A XOR2X1_32/B gnd XOR2X1_32/Y vdd XOR2X1
XXOR2X1_43 XOR2X1_43/A XOR2X1_43/B gnd XOR2X1_43/Y vdd XOR2X1
XXOR2X1_21 XOR2X1_21/A XOR2X1_21/B gnd XOR2X1_21/Y vdd XOR2X1
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B gnd XOR2X1_10/Y vdd XOR2X1
XNAND2X1_393 INVX1_312/A XOR2X1_27/Y gnd NAND3X1_403/B vdd NAND2X1
XNAND2X1_382 NAND3X1_350/C NAND3X1_350/Y gnd INVX1_322/A vdd NAND2X1
XNAND2X1_360 OR2X2_35/B OR2X2_41/A gnd AOI22X1_50/B vdd NAND2X1
XNAND2X1_371 INVX1_303/A OAI21X1_418/B gnd AOI22X1_48/B vdd NAND2X1
XINVX1_204 INVX1_204/A gnd INVX1_204/Y vdd INVX1
XINVX1_226 cos_gamma[11] gnd INVX1_226/Y vdd INVX1
XINVX1_259 cos_gamma[12] gnd INVX1_259/Y vdd INVX1
XOAI21X1_184 INVX1_28/Y INVX1_177/Y INVX1_152/A gnd OAI21X1_185/C vdd OAI21X1
XOAI21X1_151 AOI22X1_19/Y AOI22X1_20/Y AOI21X1_84/C gnd AOI21X1_70/B vdd OAI21X1
XOAI21X1_162 NOR3X1_17/B NOR3X1_17/C NOR3X1_17/A gnd AOI21X1_80/A vdd OAI21X1
XOAI21X1_195 AOI21X1_96/Y AOI21X1_97/Y AOI21X1_95/Y gnd OAI21X1_195/Y vdd OAI21X1
XOAI21X1_173 OAI21X1_173/A INVX1_171/Y AOI21X1_74/B gnd OR2X2_20/A vdd OAI21X1
XAOI22X1_5 BUFX2_3/Y vertices[5] BUFX2_16/Y vertices[4] gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_140 AOI21X1_60/Y AOI21X1_61/Y INVX1_150/Y gnd OAI21X1_140/Y vdd OAI21X1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XNAND2X1_59 XOR2X1_5/B XOR2X1_5/A gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_48 dy[4] dx[4] gnd INVX1_56/A vdd NAND2X1
XNAND2X1_15 OR2X2_4/B OR2X2_4/A gnd OAI21X1_13/C vdd NAND2X1
XNAND2X1_37 vertices[1] cos_alpha[4] gnd NOR2X1_46/A vdd NAND2X1
XNAND2X1_26 BUFX2_8/Y INVX1_43/A gnd INVX1_67/A vdd NAND2X1
XNAND2X1_190 AND2X2_46/B AND2X2_46/A gnd NAND3X1_211/A vdd NAND2X1
XAOI22X1_57 AOI22X1_57/A AOI22X1_57/B AOI22X1_57/C AOI22X1_57/D gnd AOI22X1_57/Y vdd
+ AOI22X1
XAOI21X1_208 OAI21X1_401/Y OAI21X1_431/C INVX1_315/Y gnd NOR3X1_41/B vdd AOI21X1
XAOI22X1_46 AOI22X1_46/A AOI22X1_46/B INVX1_340/A AOI22X1_46/D gnd AOI22X1_46/Y vdd
+ AOI22X1
XAOI21X1_219 AOI22X1_45/B cos_gamma[3] INVX1_342/A gnd INVX1_343/A vdd AOI21X1
XAOI22X1_35 AND2X2_67/A AOI22X1_35/B INVX1_295/A AOI22X1_35/D gnd AOI22X1_35/Y vdd
+ AOI22X1
XAOI22X1_13 NAND3X1_75/Y AOI22X1_13/B NAND3X1_77/A NAND3X1_77/C gnd NOR3X1_14/B vdd
+ AOI22X1
XAOI22X1_24 AND2X2_31/Y AND2X2_43/Y INVX1_154/Y AOI22X1_24/D gnd AOI22X1_24/Y vdd
+ AOI22X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XFILL_23_1_2 gnd vdd FILL
XOAI22X1_8 OAI22X1_8/A OAI22X1_8/B OAI22X1_8/C OAI22X1_8/D gnd OAI22X1_8/Y vdd OAI22X1
XFILL_6_2_2 gnd vdd FILL
XFILL_14_1_2 gnd vdd FILL
XAOI21X1_90 AOI21X1_90/A INVX1_212/A XNOR2X1_28/Y gnd AOI21X1_90/Y vdd AOI21X1
XFILL_19_1 gnd vdd FILL
XAND2X2_104 XNOR2X1_63/Y NOR2X1_183/A gnd NOR2X1_184/B vdd AND2X2
XNAND3X1_521 OAI21X1_482/Y NAND3X1_521/B NAND3X1_521/C gnd NAND3X1_521/Y vdd NAND3X1
XNAND3X1_532 NAND3X1_532/A NAND3X1_532/B NAND3X1_532/C gnd NAND3X1_535/A vdd NAND3X1
XNAND3X1_510 NAND3X1_510/A NAND3X1_510/B XOR2X1_43/Y gnd NAND3X1_533/B vdd NAND3X1
XNAND3X1_543 OAI21X1_511/Y NAND3X1_543/B OAI21X1_514/Y gnd NAND3X1_545/B vdd NAND3X1
XNOR2X1_200 NOR2X1_200/A NOR2X1_200/B gnd NOR3X1_48/C vdd NOR2X1
XFILL_28_0_2 gnd vdd FILL
XFILL_3_0_2 gnd vdd FILL
XFILL_19_0_2 gnd vdd FILL
XNAND3X1_384 AND2X2_93/B AOI22X1_42/D AND2X2_81/Y gnd AND2X2_93/A vdd NAND3X1
XNAND3X1_362 NOR3X1_35/A OAI21X1_347/Y NAND3X1_362/C gnd NAND3X1_362/Y vdd NAND3X1
XNAND3X1_351 OAI21X1_334/Y INVX1_284/Y OR2X2_33/Y gnd OAI21X1_386/C vdd NAND3X1
XNAND3X1_340 INVX1_269/A AND2X2_84/B NAND3X1_340/C gnd AND2X2_84/A vdd NAND3X1
XNAND3X1_373 INVX1_294/Y AND2X2_89/A NAND3X1_373/C gnd NAND3X1_378/B vdd NAND3X1
XOR2X2_38 OR2X2_38/A OR2X2_38/B gnd OR2X2_38/Y vdd OR2X2
XOR2X2_49 OR2X2_49/A OR2X2_49/B gnd OR2X2_49/Y vdd OR2X2
XNAND3X1_395 INVX1_258/Y NAND3X1_395/B OAI21X1_365/Y gnd NAND3X1_396/C vdd NAND3X1
XOR2X2_27 OR2X2_27/A OR2X2_27/B gnd OR2X2_27/Y vdd OR2X2
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd OR2X2_16/Y vdd OR2X2
XOAI21X1_514 OAI21X1_514/A NOR3X1_51/Y XNOR2X1_84/Y gnd OAI21X1_514/Y vdd OAI21X1
XOAI21X1_503 NOR3X1_45/A NOR3X1_45/B NOR3X1_45/C gnd OAI21X1_503/Y vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XNAND2X1_520 XOR2X1_48/Y XOR2X1_49/Y gnd AOI22X1_58/A vdd NAND2X1
XNAND2X1_542 AOI22X1_59/C AOI22X1_59/D gnd NOR2X1_200/B vdd NAND2X1
XNAND2X1_531 OAI21X1_499/Y OAI21X1_500/Y gnd NOR2X1_198/B vdd NAND2X1
XFILL_12_2_0 gnd vdd FILL
XNAND3X1_192 OAI21X1_196/C NAND3X1_194/B NAND3X1_194/A gnd INVX1_201/A vdd NAND3X1
XNAND3X1_170 NOR2X1_93/Y OAI21X1_171/Y OR2X2_19/Y gnd AND2X2_40/B vdd NAND3X1
XNAND3X1_181 AOI21X1_90/A INVX1_212/A XNOR2X1_28/Y gnd NAND3X1_185/B vdd NAND3X1
XOAI21X1_388 OAI21X1_388/A OAI21X1_388/B INVX1_313/A gnd OAI21X1_388/Y vdd OAI21X1
XOAI21X1_399 NOR3X1_38/B NOR3X1_38/C NOR3X1_38/A gnd OAI21X1_399/Y vdd OAI21X1
XOAI21X1_344 NOR3X1_30/A NOR3X1_30/C NOR3X1_30/B gnd OAI21X1_344/Y vdd OAI21X1
XOAI21X1_333 OAI21X1_333/A OAI21X1_442/A OAI21X1_333/C gnd OR2X2_33/A vdd OAI21X1
XOAI21X1_355 INVX1_7/Y NOR2X1_196/B OAI21X1_355/C gnd OAI21X1_355/Y vdd OAI21X1
XOAI21X1_322 NOR2X1_137/Y NOR3X1_25/C XOR2X1_22/Y gnd AND2X2_87/B vdd OAI21X1
XOAI21X1_311 OAI21X1_311/A OAI21X1_314/C AND2X2_60/A gnd INVX1_260/A vdd OAI21X1
XOAI21X1_377 INVX1_22/Y NOR2X1_197/B OAI21X1_377/C gnd AND2X2_88/B vdd OAI21X1
XOAI21X1_300 OAI21X1_301/A NOR3X1_25/Y AND2X2_65/Y gnd AOI22X1_33/D vdd OAI21X1
XOAI21X1_366 AOI22X1_38/Y XNOR2X1_37/A OAI21X1_366/C gnd NOR2X1_152/B vdd OAI21X1
XXOR2X1_44 XOR2X1_44/A XOR2X1_44/B gnd XOR2X1_44/Y vdd XOR2X1
XNAND2X1_361 AND2X2_93/B AND2X2_93/A gnd OAI21X1_414/C vdd NAND2X1
XXOR2X1_33 XOR2X1_33/A XOR2X1_33/B gnd XOR2X1_33/Y vdd XOR2X1
XNAND2X1_372 AOI22X1_48/A AOI22X1_48/B gnd NAND3X1_442/A vdd NAND2X1
XNAND2X1_350 AND2X2_79/Y OAI21X1_458/A gnd NAND2X1_351/A vdd NAND2X1
XXOR2X1_22 XOR2X1_22/A XOR2X1_22/B gnd XOR2X1_22/Y vdd XOR2X1
XXOR2X1_11 XOR2X1_11/A XOR2X1_11/B gnd XOR2X1_11/Y vdd XOR2X1
XNAND2X1_394 NAND3X1_405/Y NAND3X1_407/Y gnd NOR3X1_40/A vdd NAND2X1
XNAND2X1_383 NAND3X1_346/B INVX1_280/A gnd INVX1_314/A vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 NOR2X1_16/Y OAI21X1_7/C OR2X2_3/Y gnd AND2X2_7/A vdd NAND3X1
XFILL_26_1_0 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 INVX1_22/Y OAI22X1_8/D OAI21X1_92/B gnd OAI21X1_131/C vdd OAI21X1
XINVX1_227 cos_gamma[9] gnd OAI22X1_8/C vdd INVX1
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XOAI21X1_141 NAND3X1_77/B AOI21X1_62/Y NAND3X1_78/A gnd AOI21X1_85/C vdd OAI21X1
XOAI21X1_152 AOI22X1_19/Y AOI22X1_20/Y AOI21X1_67/Y gnd AOI21X1_95/B vdd OAI21X1
XOAI21X1_163 NOR3X1_19/B NOR3X1_19/C NOR3X1_19/A gnd AOI21X1_81/A vdd OAI21X1
XOAI21X1_196 AOI21X1_96/Y AOI21X1_97/Y OAI21X1_196/C gnd OAI21X1_196/Y vdd OAI21X1
XAOI22X1_6 INVX1_1/A vertices[6] INVX1_10/A vertices[5] gnd INVX1_101/A vdd AOI22X1
XOAI21X1_174 NOR2X1_94/Y AND2X2_41/Y INVX1_172/Y gnd AND2X2_46/A vdd OAI21X1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XOAI21X1_185 OAI22X1_7/A OAI22X1_7/B OAI21X1_185/C gnd OAI22X1_7/D vdd OAI21X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XNAND2X1_27 dy[3] dx[3] gnd INVX1_33/A vdd NAND2X1
XNAND2X1_49 OR2X2_7/B OR2X2_7/A gnd NAND2X1_50/A vdd NAND2X1
XNAND2X1_16 OAI21X1_13/C OR2X2_4/Y gnd XNOR2X1_3/B vdd NAND2X1
XNAND2X1_191 AND2X2_57/B OAI21X1_203/Y gnd OAI21X1_207/B vdd NAND2X1
XNAND2X1_38 BUFX2_4/Y vertices[3] gnd INVX1_52/A vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_180 NAND3X1_183/Y NAND3X1_184/Y gnd AOI21X1_93/C vdd NAND2X1
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_58 AOI22X1_58/A AOI22X1_58/B AOI22X1_58/C AOI22X1_58/D gnd AOI22X1_58/Y vdd
+ AOI22X1
XAOI21X1_209 OAI21X1_402/Y NAND3X1_418/B OAI21X1_380/Y gnd OAI21X1_430/B vdd AOI21X1
XAOI22X1_47 AOI22X1_47/A AOI22X1_47/B AOI22X1_47/C AOI22X1_47/D gnd AOI22X1_47/Y vdd
+ AOI22X1
XAOI22X1_36 AOI22X1_36/A AOI22X1_36/B AOI22X1_36/C AOI22X1_36/D gnd AOI22X1_36/Y vdd
+ AOI22X1
XAOI22X1_14 INVX1_155/A OR2X2_15/Y NAND3X1_82/B NAND3X1_82/C gnd AOI22X1_14/Y vdd
+ AOI22X1
XAOI22X1_25 AND2X2_46/B AND2X2_46/A AND2X2_53/B AOI22X1_25/D gnd AOI22X1_25/Y vdd
+ AOI22X1
XNOR3X1_4 NOR3X1_4/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XXNOR2X1_80 XNOR2X1_80/A XNOR2X1_80/B gnd XNOR2X1_81/B vdd XNOR2X1
XOAI22X1_9 INVX1_28/Y OAI22X1_9/B INVX1_46/Y OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XAOI21X1_80 AOI21X1_80/A AOI21X1_80/B INVX1_137/A gnd NOR3X1_19/B vdd AOI21X1
XAOI21X1_91 AOI21X1_91/A AOI21X1_91/B XNOR2X1_27/Y gnd AOI21X1_91/Y vdd AOI21X1
XFILL_19_2 gnd vdd FILL
XAND2X2_105 AND2X2_105/A AND2X2_105/B gnd NOR2X1_192/B vdd AND2X2
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XNAND3X1_522 NAND3X1_522/A OAI21X1_495/Y XOR2X1_50/Y gnd NAND3X1_523/C vdd NAND3X1
XNAND3X1_544 NAND3X1_544/A AOI22X1_60/C AOI22X1_60/D gnd NAND3X1_545/C vdd NAND3X1
XNAND3X1_500 OAI21X1_469/Y AND2X2_103/Y AOI22X1_60/B gnd NAND3X1_504/B vdd NAND3X1
XNAND3X1_533 NAND3X1_533/A NAND3X1_533/B NAND3X1_533/C gnd NAND3X1_535/B vdd NAND3X1
XNAND3X1_511 XOR2X1_37/B NAND3X1_511/B OR2X2_56/Y gnd OAI21X1_485/C vdd NAND3X1
XNAND3X1_363 INVX1_276/Y OAI21X1_379/C OAI21X1_348/Y gnd NAND3X1_364/A vdd NAND3X1
XNAND3X1_385 NAND3X1_387/A AND2X2_93/A OAI21X1_363/C gnd AND2X2_94/B vdd NAND3X1
XNAND3X1_341 INVX1_269/Y NAND3X1_341/B NAND3X1_341/C gnd AND2X2_81/B vdd NAND3X1
XNAND3X1_374 NAND3X1_378/B AND2X2_80/Y OAI21X1_359/Y gnd NAND3X1_380/C vdd NAND3X1
XNAND3X1_352 OAI21X1_336/Y OAI21X1_386/C OR2X2_34/Y gnd AND2X2_74/B vdd NAND3X1
XNAND3X1_396 INVX1_297/Y NAND3X1_396/B NAND3X1_396/C gnd AOI22X1_44/B vdd NAND3X1
XNAND3X1_330 OAI21X1_304/C NAND3X1_330/B NAND3X1_330/C gnd NAND3X1_331/B vdd NAND3X1
XOR2X2_39 OR2X2_39/A OR2X2_39/B gnd OR2X2_39/Y vdd OR2X2
XOR2X2_28 OR2X2_28/A OR2X2_28/B gnd OR2X2_28/Y vdd OR2X2
XOR2X2_17 OR2X2_17/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XOAI21X1_515 OAI21X1_518/A NOR3X1_52/Y OAI21X1_515/C gnd OAI21X1_515/Y vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_504 OAI21X1_504/A NOR2X1_198/Y INVX1_378/A gnd OAI21X1_504/Y vdd OAI21X1
XNAND2X1_521 OAI21X1_492/Y NAND3X1_515/Y gnd INVX1_376/A vdd NAND2X1
XNAND2X1_543 NAND3X1_546/Y OAI21X1_515/Y gnd OAI21X1_517/C vdd NAND2X1
XNAND2X1_532 cos_gamma[3] NAND3X1_369/C gnd NOR2X1_198/A vdd NAND2X1
XNAND2X1_510 cos_alpha[3] vertices[12] gnd XOR2X1_47/B vdd NAND2X1
XFILL_12_2_1 gnd vdd FILL
XNAND3X1_160 XOR2X1_10/Y AOI21X1_74/A AOI21X1_74/B gnd NAND3X1_163/B vdd NAND3X1
XNAND3X1_193 INVX1_201/A OAI21X1_195/Y INVX1_173/Y gnd INVX1_216/A vdd NAND3X1
XNAND3X1_171 INVX1_172/A OAI21X1_213/C OR2X2_20/Y gnd AND2X2_46/B vdd NAND3X1
XNAND3X1_182 NAND3X1_185/A OAI21X1_192/C NAND3X1_185/B gnd INVX1_213/A vdd NAND3X1
XOAI21X1_312 INVX1_259/Y INVX1_9/Y INVX1_260/Y gnd AND2X2_66/B vdd OAI21X1
XOAI21X1_323 NOR2X1_137/Y NOR3X1_25/C XNOR2X1_38/Y gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_301 OAI21X1_301/A NOR3X1_25/Y OAI21X1_301/C gnd AOI22X1_34/D vdd OAI21X1
XOAI21X1_389 NOR3X1_31/A NOR3X1_31/B OAI21X1_389/C gnd OAI21X1_389/Y vdd OAI21X1
XOAI21X1_345 NOR3X1_31/A NOR3X1_31/C NOR3X1_31/B gnd OAI21X1_345/Y vdd OAI21X1
XOAI21X1_378 NOR2X1_137/B NOR2X1_173/A AND2X2_89/A gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_334 INVX1_50/Y NOR2X1_86/B OR2X2_33/A gnd OAI21X1_334/Y vdd OAI21X1
XOAI21X1_356 INVX1_7/Y NOR2X1_196/B OAI21X1_356/C gnd OAI21X1_356/Y vdd OAI21X1
XOAI21X1_367 INVX1_298/Y INVX1_9/Y OAI21X1_475/A gnd OAI21X1_368/C vdd OAI21X1
XNAND2X1_384 vertices[1] cos_alpha[12] gnd OAI21X1_491/A vdd NAND2X1
XXOR2X1_23 XOR2X1_23/A XOR2X1_23/B gnd XOR2X1_23/Y vdd XOR2X1
XXOR2X1_45 XOR2X1_45/A XOR2X1_45/B gnd XOR2X1_45/Y vdd XOR2X1
XXOR2X1_34 XOR2X1_34/A XOR2X1_34/B gnd XOR2X1_35/A vdd XOR2X1
XNAND2X1_373 AND2X2_92/B AND2X2_92/A gnd OAI21X1_411/C vdd NAND2X1
XNAND2X1_395 vertices[5] cos_alpha[8] gnd OR2X2_39/B vdd NAND2X1
XNAND2X1_351 NAND2X1_351/A NAND2X1_351/B gnd NAND3X1_369/C vdd NAND2X1
XNAND2X1_340 cos_alpha[3] vertices[9] gnd AND2X2_75/B vdd NAND2X1
XNAND2X1_362 cos_gamma[9] AND2X2_13/Y gnd OAI21X1_476/A vdd NAND2X1
XXOR2X1_12 XOR2X1_12/A XOR2X1_12/B gnd XOR2X1_12/Y vdd XOR2X1
XNAND3X1_2 BUFX2_7/Y NOR2X1_7/Y INVX1_18/A gnd NAND3X1_2/Y vdd NAND3X1
XFILL_26_1_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_120 NOR3X1_10/B NOR3X1_9/Y NOR3X1_10/A gnd AOI21X1_53/A vdd OAI21X1
XOAI21X1_153 AOI21X1_69/Y AOI21X1_70/Y AOI21X1_68/Y gnd OAI21X1_153/Y vdd OAI21X1
XOAI21X1_164 NOR3X1_17/A NOR3X1_17/B AOI21X1_78/B gnd INVX1_191/A vdd OAI21X1
XAOI22X1_7 INVX1_102/Y INVX1_103/Y INVX1_74/Y AOI22X1_7/D gnd NOR3X1_4/A vdd AOI22X1
XOAI21X1_131 OR2X2_18/B OR2X2_19/B OAI21X1_131/C gnd OR2X2_16/A vdd OAI21X1
XOAI21X1_142 INVX1_50/Y INVX1_46/Y OAI22X1_7/A gnd AOI22X1_23/D vdd OAI21X1
XINVX1_228 INVX1_228/A gnd INVX1_228/Y vdd INVX1
XINVX1_206 OAI22X1_7/Y gnd INVX1_206/Y vdd INVX1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XOAI21X1_197 INVX1_157/Y NOR2X1_89/A INVX1_158/A gnd XOR2X1_11/B vdd OAI21X1
XOAI21X1_175 INVX1_155/A AOI21X1_84/Y INVX1_183/A gnd OAI21X1_196/C vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_186 INVX1_154/A NOR2X1_97/Y AOI22X1_17/D gnd OAI21X1_189/C vdd OAI21X1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XNAND2X1_17 AND2X2_4/Y XOR2X1_3/Y gnd INVX1_21/A vdd NAND2X1
XNAND2X1_28 OR2X2_5/B OR2X2_5/A gnd NAND2X1_29/A vdd NAND2X1
XNAND2X1_192 NAND3X1_275/A OAI21X1_205/Y gnd NAND2X1_193/B vdd NAND2X1
XNAND2X1_39 INVX1_10/A vertices[4] gnd OAI21X1_43/C vdd NAND2X1
XNAND2X1_181 NAND3X1_199/Y OAI21X1_219/C gnd NOR2X1_107/B vdd NAND2X1
XNAND2X1_170 OR2X2_21/B OR2X2_21/A gnd INVX1_202/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_59 OR2X2_55/Y AOI22X1_59/B AOI22X1_59/C AOI22X1_59/D gnd NOR3X1_48/A vdd
+ AOI22X1
XAOI22X1_48 AOI22X1_48/A AOI22X1_48/B AOI22X1_48/C AOI22X1_48/D gnd AOI22X1_48/Y vdd
+ AOI22X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_6/C vdd NOR3X1
XAOI22X1_15 cos_gamma[2] NAND2X1_70/Y AOI22X1_15/C AND2X2_36/B gnd NOR3X1_5/B vdd
+ AOI22X1
XAOI22X1_26 OR2X2_17/Y AND2X2_47/B AND2X2_56/B AOI22X1_26/D gnd AOI22X1_26/Y vdd AOI22X1
XAOI22X1_37 AOI22X1_37/A OR2X2_27/Y AOI22X1_37/C AOI22X1_37/D gnd AOI22X1_37/Y vdd
+ AOI22X1
XXNOR2X1_81 XNOR2X1_81/A XNOR2X1_81/B gnd XOR2X1_51/A vdd XNOR2X1
XXNOR2X1_70 XNOR2X1_70/A XNOR2X1_70/B gnd XNOR2X1_71/A vdd XNOR2X1
XAOI21X1_70 AOI21X1_70/A AOI21X1_70/B INVX1_155/A gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_81 AOI21X1_81/A XNOR2X1_23/B NOR3X1_19/Y gnd XOR2X1_12/B vdd AOI21X1
XAOI21X1_92 AOI21X1_92/A INVX1_213/A AOI21X1_92/C gnd AOI21X1_92/Y vdd AOI21X1
XAND2X2_106 XOR2X1_46/A XOR2X1_46/B gnd AND2X2_106/Y vdd AND2X2
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd XOR2X1_3/A vdd XOR2X1
XFILL_6_0_1 gnd vdd FILL
XNAND3X1_545 INVX1_384/Y NAND3X1_545/B NAND3X1_545/C gnd NAND3X1_547/A vdd NAND3X1
XNAND3X1_523 NAND3X1_523/A NAND3X1_523/B NAND3X1_523/C gnd NAND3X1_523/Y vdd NAND3X1
XNAND3X1_501 OR2X2_35/Y NAND3X1_504/B OAI21X1_471/Y gnd NAND3X1_502/B vdd NAND3X1
XNAND3X1_512 OAI21X1_445/Y OR2X2_51/Y XNOR2X1_50/A gnd AND2X2_105/B vdd NAND3X1
XNAND3X1_534 NAND3X1_534/A INVX1_379/A OR2X2_59/Y gnd AND2X2_109/B vdd NAND3X1
XFILL_24_1 gnd vdd FILL
XNAND3X1_364 NAND3X1_364/A OAI21X1_350/Y INVX1_290/Y gnd NAND3X1_423/A vdd NAND3X1
XNAND3X1_386 AND2X2_94/B AOI22X1_43/D INVX1_264/Y gnd AND2X2_94/A vdd NAND3X1
XNAND3X1_353 INVX1_285/A OAI21X1_339/Y INVX1_286/Y gnd AND2X2_77/A vdd NAND3X1
XNAND3X1_342 INVX1_272/Y NAND3X1_375/B AND2X2_87/B gnd NAND3X1_342/Y vdd NAND3X1
XNAND3X1_375 INVX1_272/A NAND3X1_375/B AND2X2_87/B gnd AND2X2_87/A vdd NAND3X1
XNAND3X1_397 cos_gamma[9] NOR2X1_131/Y AND2X2_13/Y gnd AND2X2_97/B vdd NAND3X1
XNAND3X1_320 AOI22X1_34/C NAND3X1_320/B AOI22X1_34/D gnd NAND3X1_326/A vdd NAND3X1
XNAND3X1_331 INVX1_225/A NAND3X1_331/B OAI21X1_305/Y gnd NAND3X1_334/C vdd NAND3X1
XOR2X2_29 OR2X2_29/A OR2X2_29/B gnd OR2X2_29/Y vdd OR2X2
XOR2X2_18 OR2X2_19/B OR2X2_18/B gnd OR2X2_18/Y vdd OR2X2
XFILL_21_2_2 gnd vdd FILL
XOAI21X1_505 INVX1_333/Y XNOR2X1_47/A OR2X2_46/Y gnd INVX1_379/A vdd OAI21X1
XOAI21X1_516 NOR3X1_52/B NOR3X1_52/C NOR3X1_52/A gnd OAI21X1_516/Y vdd OAI21X1
XNAND2X1_522 AOI22X1_58/D AOI22X1_58/C gnd NAND3X1_517/A vdd NAND2X1
XNAND2X1_544 NOR2X1_178/A NOR2X1_178/B gnd NAND3X1_548/C vdd NAND2X1
XNAND2X1_500 NAND3X1_533/B NAND3X1_533/A gnd NAND3X1_532/C vdd NAND2X1
XNAND2X1_533 NAND3X1_532/B NAND3X1_532/A gnd NAND3X1_533/C vdd NAND2X1
XNAND2X1_511 INVX1_15/A vertices[13] gnd XNOR2X1_71/B vdd NAND2X1
XFILL_12_2_2 gnd vdd FILL
XAOI21X1_190 NAND3X1_327/A AOI22X1_35/D INVX1_295/Y gnd OAI21X1_362/C vdd AOI21X1
XNAND3X1_150 NAND3X1_99/C NAND3X1_200/A NAND3X1_150/C gnd NAND3X1_155/B vdd NAND3X1
XNAND3X1_161 NAND3X1_163/B OAI21X1_157/Y INVX1_161/Y gnd AOI21X1_76/B vdd NAND3X1
XNAND3X1_194 NAND3X1_194/A NAND3X1_194/B AOI21X1_95/Y gnd NAND3X1_198/A vdd NAND3X1
XNAND3X1_172 OAI21X1_180/Y INVX1_176/Y OR2X2_22/Y gnd NAND3X1_183/B vdd NAND3X1
XNAND3X1_183 INVX1_175/A NAND3X1_183/B OAI21X1_181/Y gnd NAND3X1_183/Y vdd NAND3X1
XOAI21X1_324 INVX1_29/Y NOR2X1_95/B XOR2X1_23/A gnd OAI21X1_325/C vdd OAI21X1
XOAI21X1_346 NOR3X1_32/B NOR3X1_32/C NOR3X1_32/A gnd OAI21X1_346/Y vdd OAI21X1
XOAI21X1_335 NOR3X1_26/Y OAI21X1_386/B NOR2X1_143/Y gnd AND2X2_74/A vdd OAI21X1
XOAI21X1_313 INVX1_232/Y NOR2X1_116/A INVX1_231/A gnd INVX1_269/A vdd OAI21X1
XOAI21X1_302 AOI22X1_33/Y AOI22X1_34/Y OAI21X1_302/C gnd AOI22X1_36/D vdd OAI21X1
XOAI21X1_357 INVX1_250/Y NOR2X1_128/A INVX1_251/A gnd XOR2X1_24/B vdd OAI21X1
XOAI21X1_379 INVX1_276/A OAI21X1_379/B OAI21X1_379/C gnd OAI21X1_379/Y vdd OAI21X1
XOAI21X1_368 NOR2X1_163/A INVX1_299/Y OAI21X1_368/C gnd XOR2X1_25/B vdd OAI21X1
XNAND2X1_385 vertices[1] cos_alpha[13] gnd OR2X2_48/B vdd NAND2X1
XXOR2X1_35 XOR2X1_35/A XOR2X1_35/B gnd OR2X2_50/A vdd XOR2X1
XXOR2X1_46 XOR2X1_46/A XOR2X1_46/B gnd XOR2X1_46/Y vdd XOR2X1
XXOR2X1_24 XOR2X1_24/A XOR2X1_24/B gnd XOR2X1_24/Y vdd XOR2X1
XNAND2X1_341 AND2X2_77/B AND2X2_77/A gnd NOR3X1_29/B vdd NAND2X1
XNAND2X1_396 cos_alpha[6] vertices[7] gnd OAI21X1_484/A vdd NAND2X1
XNAND2X1_352 OAI21X1_406/A OAI21X1_458/A gnd NAND2X1_353/A vdd NAND2X1
XNAND2X1_330 XOR2X1_18/A INVX1_275/Y gnd INVX1_276/A vdd NAND2X1
XNAND2X1_374 cos_gamma[5] NAND3X1_457/B gnd XOR2X1_26/B vdd NAND2X1
XXOR2X1_13 XOR2X1_13/A XOR2X1_13/B gnd XOR2X1_13/Y vdd XOR2X1
XNAND2X1_363 cos_gamma[6] NAND2X1_536/B gnd NOR2X1_169/A vdd NAND2X1
XNAND3X1_3 INVX1_17/A INVX1_31/A NAND3X1_3/C gnd NAND3X1_3/Y vdd NAND3X1
XFILL_26_1_2 gnd vdd FILL
XFILL_1_1_2 gnd vdd FILL
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XOAI21X1_121 AOI21X1_53/Y NOR3X1_11/Y OR2X2_12/Y gnd AOI22X1_16/D vdd OAI21X1
XOAI21X1_110 INVX1_8/Y INVX1_124/Y AOI21X1_43/Y gnd AOI21X1_45/A vdd OAI21X1
XOAI21X1_154 AOI21X1_69/Y AOI21X1_70/Y OAI21X1_154/C gnd AOI21X1_83/A vdd OAI21X1
XAOI22X1_8 BUFX2_12/Y vertices[4] INVX1_101/Y AOI22X1_8/D gnd NOR3X1_4/C vdd AOI22X1
XOAI21X1_165 INVX1_140/Y AOI21X1_75/Y INVX1_162/A gnd INVX1_190/A vdd OAI21X1
XOAI21X1_198 NOR3X1_20/B NOR3X1_20/C NOR3X1_20/A gnd OAI21X1_198/Y vdd OAI21X1
XOAI21X1_132 INVX1_65/Y INVX1_43/Y OR2X2_16/A gnd AND2X2_35/B vdd OAI21X1
XOAI21X1_176 OAI21X1_176/A AOI21X1_85/Y INVX1_182/A gnd OAI21X1_193/C vdd OAI21X1
XOAI21X1_143 NOR2X1_76/B INVX1_152/A AOI22X1_23/D gnd XNOR2X1_21/A vdd OAI21X1
XOAI21X1_187 INVX1_10/Y OAI22X1_6/D AND2X2_44/Y gnd AOI21X1_88/A vdd OAI21X1
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XINVX1_218 dz[10] gnd INVX1_218/Y vdd INVX1
XFILL_9_2_2 gnd vdd FILL
XFILL_17_1_2 gnd vdd FILL
XNAND2X1_18 XOR2X1_2/B XOR2X1_2/A gnd NAND2X1_20/A vdd NAND2X1
XNAND2X1_29 NAND2X1_29/A OR2X2_5/Y gnd OR2X2_6/A vdd NAND2X1
XNAND2X1_160 AOI22X1_22/C AOI21X1_75/A gnd INVX1_189/A vdd NAND2X1
XNAND2X1_193 NAND3X1_169/Y NAND2X1_193/B gnd NAND2X1_194/B vdd NAND2X1
XNAND2X1_171 INVX1_202/A OR2X2_21/Y gnd AOI21X1_97/C vdd NAND2X1
XNAND2X1_182 NOR2X1_107/B NAND2X1_185/B gnd AOI21X1_98/A vdd NAND2X1
XAOI22X1_49 AOI22X1_49/A AOI22X1_49/B AOI22X1_49/C AOI22X1_49/D gnd AOI22X1_49/Y vdd
+ AOI22X1
XAOI22X1_27 INVX1_208/Y NOR2X1_97/B INVX1_178/Y OAI22X1_6/Y gnd INVX1_211/A vdd AOI22X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_7/C vdd NOR3X1
XAOI22X1_16 INVX1_112/Y NOR2X1_66/Y NOR3X1_19/A AOI22X1_16/D gnd NOR2X1_81/A vdd AOI22X1
XAOI22X1_38 AOI22X1_38/A INVX1_257/Y INVX1_297/A AOI22X1_38/D gnd AOI22X1_38/Y vdd
+ AOI22X1
XXNOR2X1_82 INVX1_366/A OR2X2_54/B gnd NOR3X1_50/B vdd XNOR2X1
XXNOR2X1_60 XOR2X1_42/Y dx[15] gnd XOR2X1_43/B vdd XNOR2X1
XXNOR2X1_71 XNOR2X1_71/A XNOR2X1_71/B gnd XNOR2X1_72/A vdd XNOR2X1
XAOI21X1_71 NAND3X1_93/C NAND3X1_93/A INVX1_125/A gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_82 AOI21X1_82/A AOI21X1_82/B INVX1_8/Y gnd INVX1_171/A vdd AOI21X1
XAOI21X1_93 AOI21X1_93/A AOI21X1_93/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XAOI21X1_60 AOI21X1_60/A AOI21X1_60/B NOR2X1_86/Y gnd AOI21X1_60/Y vdd AOI21X1
XAND2X2_107 OR2X2_58/A OR2X2_58/B gnd OAI22X1_13/D vdd AND2X2
XFILL_6_0_2 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd XOR2X1_3/Y vdd XOR2X1
XNAND3X1_546 NAND3X1_547/A OAI21X1_518/C OAI21X1_516/Y gnd NAND3X1_546/Y vdd NAND3X1
XNAND3X1_502 NAND3X1_502/A NAND3X1_502/B AND2X2_96/Y gnd AOI22X1_56/A vdd NAND3X1
XNAND3X1_535 NAND3X1_535/A NAND3X1_535/B AND2X2_109/Y gnd NAND3X1_536/B vdd NAND3X1
XNAND3X1_524 NAND3X1_524/A OR2X2_58/Y NAND3X1_524/C gnd AND2X2_108/A vdd NAND3X1
XNAND3X1_513 OR2X2_57/Y OR2X2_52/Y XOR2X1_46/Y gnd NAND3X1_513/Y vdd NAND3X1
XFILL_24_2 gnd vdd FILL
XFILL_17_1 gnd vdd FILL
XFILL_24_2_0 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XNAND3X1_310 INVX1_239/A OAI21X1_296/C AOI22X1_41/D gnd NAND3X1_311/C vdd NAND3X1
XNAND3X1_321 INVX1_270/A NAND3X1_321/B AOI22X1_33/D gnd NAND3X1_326/B vdd NAND3X1
XNAND3X1_332 NAND3X1_334/B NAND3X1_334/C OAI21X1_307/C gnd INVX1_297/A vdd NAND3X1
XNAND3X1_354 INVX1_287/Y INVX1_288/Y OAI21X1_395/C gnd NAND3X1_412/B vdd NAND3X1
XNAND3X1_387 NAND3X1_387/A OAI21X1_362/C AND2X2_93/A gnd NAND3X1_388/B vdd NAND3X1
XNAND3X1_365 INVX1_291/Y OAI21X1_352/Y NAND3X1_423/A gnd INVX1_359/A vdd NAND3X1
XNAND3X1_398 cos_gamma[11] INVX1_18/A INVX1_304/A gnd AND2X2_97/A vdd NAND3X1
XNAND3X1_376 INVX1_272/Y NAND3X1_376/B OAI21X1_323/Y gnd NAND3X1_376/Y vdd NAND3X1
XNAND3X1_343 INVX1_272/A NAND3X1_376/B OAI21X1_323/Y gnd NAND3X1_343/Y vdd NAND3X1
XOR2X2_19 OR2X2_19/A OR2X2_19/B gnd OR2X2_19/Y vdd OR2X2
XOAI21X1_517 INVX1_386/A NOR2X1_179/A OAI21X1_517/C gnd OAI21X1_517/Y vdd OAI21X1
XOAI21X1_506 INVX1_336/Y INVX1_337/Y INVX1_338/Y gnd XNOR2X1_78/A vdd OAI21X1
XNAND2X1_523 NAND3X1_522/A OAI21X1_495/Y gnd NAND2X1_525/B vdd NAND2X1
XNAND2X1_545 NAND3X1_547/Y OAI21X1_518/Y gnd NAND3X1_548/B vdd NAND2X1
XNAND2X1_501 OR2X2_56/B OR2X2_56/A gnd NAND3X1_511/B vdd NAND2X1
XNAND2X1_534 cos_gamma[9] NOR2X1_73/Y gnd XNOR2X1_78/B vdd NAND2X1
XNAND2X1_512 BUFX2_4/Y vertices[15] gnd XNOR2X1_70/B vdd NAND2X1
XAOI21X1_180 OAI21X1_346/Y OAI21X1_380/C INVX1_282/Y gnd NOR3X1_35/B vdd AOI21X1
XAOI21X1_191 OAI21X1_360/Y NAND3X1_382/A NAND3X1_382/B gnd OAI21X1_363/B vdd AOI21X1
XNAND3X1_140 INVX1_155/Y INVX1_183/A AOI21X1_95/B gnd NAND3X1_144/B vdd NAND3X1
XNAND3X1_151 AOI21X1_56/Y NAND3X1_151/B NAND3X1_151/C gnd NAND3X1_155/C vdd NAND3X1
XNAND3X1_162 AOI21X1_76/B AOI21X1_76/C AOI21X1_76/A gnd AOI21X1_75/B vdd NAND3X1
XNAND3X1_184 INVX1_175/Y NAND3X1_184/B OAI21X1_182/Y gnd NAND3X1_184/Y vdd NAND3X1
XNAND3X1_173 INVX1_175/Y NAND3X1_183/B OAI21X1_181/Y gnd NAND3X1_173/Y vdd NAND3X1
XNAND3X1_195 INVX1_173/A NAND3X1_198/A OAI21X1_196/Y gnd NAND3X1_200/B vdd NAND3X1
XOAI21X1_325 OAI21X1_325/A OAI21X1_325/B OAI21X1_325/C gnd OAI21X1_326/C vdd OAI21X1
XOAI21X1_347 NOR3X1_33/B NOR3X1_33/C NOR3X1_33/A gnd OAI21X1_347/Y vdd OAI21X1
XOAI21X1_369 NOR2X1_163/A INVX1_260/Y INVX1_300/Y gnd AND2X2_83/B vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_358 OAI21X1_359/A OAI21X1_359/B INVX1_294/Y gnd OAI21X1_358/Y vdd OAI21X1
XOAI21X1_336 NOR3X1_26/B NOR3X1_26/C NOR3X1_26/A gnd OAI21X1_336/Y vdd OAI21X1
XOAI21X1_314 OAI22X1_8/C INVX1_43/Y OAI21X1_314/C gnd AND2X2_68/B vdd OAI21X1
XOAI21X1_303 AOI22X1_33/Y AOI22X1_34/Y OAI21X1_303/C gnd AOI22X1_35/D vdd OAI21X1
XXOR2X1_36 XOR2X1_36/A XOR2X1_36/B gnd XOR2X1_36/Y vdd XOR2X1
XXOR2X1_25 XOR2X1_25/A XOR2X1_25/B gnd XOR2X1_25/Y vdd XOR2X1
XNAND2X1_320 cos_gamma[5] NAND2X1_536/B gnd XOR2X1_22/B vdd NAND2X1
XXOR2X1_14 XOR2X1_14/A XOR2X1_14/B gnd XOR2X1_14/Y vdd XOR2X1
XNAND2X1_386 vertices[2] cos_alpha[11] gnd OR2X2_38/B vdd NAND2X1
XNAND2X1_375 cos_gamma[1] NAND3X1_369/C gnd NOR2X1_173/A vdd NAND2X1
XNAND2X1_397 vertices[7] cos_alpha[7] gnd OAI21X1_443/C vdd NAND2X1
XNAND2X1_353 NAND2X1_353/A NAND3X1_429/C gnd NOR2X1_196/B vdd NAND2X1
XNAND2X1_331 INVX1_289/A NAND3X1_301/B gnd OAI21X1_349/C vdd NAND2X1
XNAND2X1_342 BUFX2_12/Y vertices[10] gnd NOR3X1_27/A vdd NAND2X1
XXOR2X1_47 OR2X2_57/B XOR2X1_47/B gnd XOR2X1_47/Y vdd XOR2X1
XNAND2X1_364 cos_gamma[7] NAND2X1_536/B gnd NOR2X1_166/B vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_4 INVX1_51/Y NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_5/A vdd NAND3X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XAOI22X1_9 AOI22X1_9/A AOI22X1_9/B AOI22X1_9/C AOI22X1_9/D gnd NOR3X1_3/A vdd AOI22X1
XOAI21X1_122 NOR3X1_11/B NOR3X1_11/C INVX1_92/Y gnd OAI21X1_122/Y vdd OAI21X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XOAI21X1_155 INVX1_130/Y NOR2X1_80/A INVX1_131/A gnd XOR2X1_10/B vdd OAI21X1
XOAI21X1_111 INVX1_8/Y INVX1_124/Y OAI21X1_173/A gnd AOI22X1_15/C vdd OAI21X1
XOAI21X1_133 OR2X2_11/A INVX1_142/Y AND2X2_36/A gnd OAI21X1_133/Y vdd OAI21X1
XOAI21X1_100 INVX1_100/A INVX1_101/A AOI22X1_8/D gnd NAND3X1_72/A vdd OAI21X1
XOAI21X1_199 OAI21X1_200/A NOR3X1_20/Y INVX1_188/Y gnd AOI22X1_25/D vdd OAI21X1
XOAI21X1_144 INVX1_29/Y INVX1_71/Y XNOR2X1_21/A gnd AOI22X1_18/B vdd OAI21X1
XOAI21X1_166 INVX1_91/Y INVX1_43/Y OAI22X1_5/B gnd OAI21X1_167/C vdd OAI21X1
XOAI21X1_177 NOR2X1_74/B INVX1_147/A OAI21X1_177/C gnd INVX1_175/A vdd OAI21X1
XOAI21X1_188 INVX1_1/Y OAI22X1_6/B AND2X2_43/Y gnd AOI21X1_88/B vdd OAI21X1
XNAND2X1_19 XOR2X1_3/B XOR2X1_3/A gnd NAND2X1_20/B vdd NAND2X1
XNAND2X1_150 cos_gamma[2] NOR2X1_73/Y gnd INVX1_160/A vdd NAND2X1
XNAND2X1_161 cos_gamma[3] NOR2X1_73/Y gnd OR2X2_19/A vdd NAND2X1
XNAND2X1_172 vertices[3] cos_alpha[7] gnd INVX1_205/A vdd NAND2X1
XNAND2X1_194 OAI21X1_308/C NAND2X1_194/B gnd XOR2X1_12/A vdd NAND2X1
XNAND2X1_183 NAND3X1_200/Y NAND3X1_201/Y gnd NAND3X1_202/C vdd NAND2X1
XAOI22X1_39 AOI22X1_39/A AOI22X1_39/B AOI22X1_39/C AOI22X1_39/D gnd AOI22X1_39/Y vdd
+ AOI22X1
XAOI22X1_17 BUFX2_11/Y vertices[6] AOI22X1_24/D AOI22X1_17/D gnd AOI22X1_17/Y vdd
+ AOI22X1
XAOI22X1_28 AND2X2_61/A AND2X2_54/B INVX1_253/A AOI22X1_28/D gnd AOI22X1_28/Y vdd
+ AOI22X1
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_8/C vdd NOR3X1
XXNOR2X1_83 NOR3X1_48/B INVX1_383/Y gnd XNOR2X1_83/Y vdd XNOR2X1
XXNOR2X1_61 XOR2X1_43/A XOR2X1_43/B gnd XNOR2X1_61/Y vdd XNOR2X1
XXNOR2X1_50 XNOR2X1_50/A XNOR2X1_50/B gnd XOR2X1_36/A vdd XNOR2X1
XXNOR2X1_72 XNOR2X1_72/A XOR2X1_47/Y gnd XOR2X1_49/A vdd XNOR2X1
XFILL_5_1 gnd vdd FILL
XAOI21X1_50 OAI21X1_83/Y INVX1_118/A INVX1_110/A gnd AOI21X1_50/Y vdd AOI21X1
XAOI21X1_72 NAND3X1_98/C NAND3X1_98/B NAND3X1_95/A gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_83 AOI21X1_83/A AOI21X1_83/B NAND3X1_96/C gnd AOI21X1_83/Y vdd AOI21X1
XOAI21X1_1 INVX1_2/Y INVX1_10/Y OAI21X1_7/A gnd OAI21X1_2/C vdd OAI21X1
XAOI21X1_94 AOI21X1_94/A AOI22X1_19/D INVX1_182/Y gnd AOI21X1_94/Y vdd AOI21X1
XAOI21X1_61 AOI21X1_61/A AOI21X1_61/B INVX1_145/Y gnd AOI21X1_61/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XAND2X2_108 AND2X2_108/A OAI22X1_13/Y gnd AND2X2_108/Y vdd AND2X2
XNAND3X1_514 INVX1_373/A OAI22X1_10/Y OAI22X1_11/Y gnd NAND3X1_516/C vdd NAND3X1
XNAND3X1_503 OR2X2_35/Y INVX1_385/A OAI21X1_470/Y gnd NAND3X1_505/B vdd NAND3X1
XXOR2X1_4 XOR2X1_4/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XNAND3X1_547 NAND3X1_547/A OAI21X1_516/Y OAI21X1_515/C gnd NAND3X1_547/Y vdd NAND3X1
XNAND3X1_536 XNOR2X1_59/Y NAND3X1_536/B OAI21X1_507/Y gnd AOI22X1_59/C vdd NAND3X1
XNAND3X1_525 OAI21X1_499/Y OAI21X1_500/Y NOR2X1_196/Y gnd NAND3X1_530/A vdd NAND3X1
XFILL_17_2 gnd vdd FILL
XINVX1_380 NOR3X1_48/A gnd INVX1_380/Y vdd INVX1
XFILL_24_2_1 gnd vdd FILL
XNAND3X1_344 OAI21X1_326/Y INVX1_278/Y NAND3X1_344/C gnd NAND3X1_346/B vdd NAND3X1
XNAND3X1_355 OAI21X1_341/Y NAND3X1_412/B OAI21X1_340/Y gnd NAND3X1_356/A vdd NAND3X1
XNAND3X1_366 BUFX2_8/Y OAI21X1_356/C NAND3X1_369/C gnd NAND3X1_368/B vdd NAND3X1
XNAND3X1_311 INVX1_7/A OAI21X1_297/Y NAND3X1_311/C gnd NOR2X1_137/B vdd NAND3X1
XNAND3X1_300 NAND3X1_301/B OAI21X1_293/C NAND3X1_301/A gnd INVX1_274/A vdd NAND3X1
XFILL_15_2_1 gnd vdd FILL
XNAND3X1_322 OAI21X1_303/C NAND3X1_326/A NAND3X1_326/B gnd AOI22X1_36/C vdd NAND3X1
XNAND3X1_333 INVX1_256/A INVX1_297/A AOI22X1_38/D gnd AOI22X1_39/C vdd NAND3X1
XNAND3X1_388 INVX1_264/A NAND3X1_388/B OAI21X1_363/Y gnd NAND3X1_391/A vdd NAND3X1
XNAND3X1_377 NAND3X1_377/A AND2X2_80/Y OAI21X1_358/Y gnd NAND3X1_379/B vdd NAND3X1
XNAND3X1_399 cos_gamma[4] NAND3X1_399/B NOR2X1_157/Y gnd AND2X2_88/A vdd NAND3X1
XOAI21X1_518 OAI21X1_518/A NOR3X1_52/Y OAI21X1_518/C gnd OAI21X1_518/Y vdd OAI21X1
XOAI21X1_507 NOR3X1_47/B NOR3X1_47/C NOR3X1_47/A gnd OAI21X1_507/Y vdd OAI21X1
XNAND2X1_502 vertices[3] cos_alpha[12] gnd XNOR2X1_63/B vdd NAND2X1
XNAND2X1_546 NAND3X1_548/Y OAI21X1_517/Y gnd NAND2X1_546/Y vdd NAND2X1
XNAND2X1_524 XOR2X1_50/Y NAND2X1_525/B gnd NAND3X1_521/B vdd NAND2X1
XNAND2X1_513 NOR2X1_191/A XOR2X1_45/Y gnd AOI22X1_57/C vdd NAND2X1
XNAND2X1_535 cos_gamma[6] NAND3X1_399/B gnd XOR2X1_51/B vdd NAND2X1
XAOI21X1_181 OAI21X1_348/Y OAI21X1_379/C INVX1_276/Y gnd NOR3X1_34/B vdd AOI21X1
XAOI21X1_192 OAI21X1_363/Y NAND3X1_388/B INVX1_264/A gnd OAI21X1_365/B vdd AOI21X1
XAOI21X1_170 OAI21X1_281/Y INVX1_244/Y NOR2X1_125/Y gnd NOR3X1_28/A vdd AOI21X1
XNAND3X1_141 NAND3X1_144/B OAI21X1_154/C NAND3X1_144/A gnd INVX1_173/A vdd NAND3X1
XNAND3X1_163 INVX1_161/A NAND3X1_163/B OAI21X1_157/Y gnd AOI22X1_22/C vdd NAND3X1
XNAND3X1_152 AOI21X1_72/Y NAND3X1_155/B NAND3X1_155/C gnd AOI21X1_82/A vdd NAND3X1
XNAND3X1_196 AOI21X1_83/Y NAND3X1_200/B INVX1_216/A gnd OAI21X1_219/C vdd NAND3X1
XNAND3X1_130 INVX1_181/A AOI22X1_18/D XNOR2X1_21/Y gnd AOI21X1_85/A vdd NAND3X1
XNAND3X1_185 NAND3X1_185/A NAND3X1_185/B AOI21X1_89/Y gnd AOI21X1_93/B vdd NAND3X1
XNAND3X1_174 OAI21X1_180/Y INVX1_176/A OR2X2_22/Y gnd NAND3X1_184/B vdd NAND3X1
XOAI21X1_326 INVX1_45/Y INVX1_241/Y OAI21X1_326/C gnd OAI21X1_326/Y vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_348 NOR3X1_35/B NOR3X1_35/C NOR3X1_35/A gnd OAI21X1_348/Y vdd OAI21X1
XOAI21X1_359 OAI21X1_359/A OAI21X1_359/B XOR2X1_24/Y gnd OAI21X1_359/Y vdd OAI21X1
XOAI21X1_315 INVX1_226/Y NOR2X1_7/B INVX1_265/Y gnd AND2X2_69/A vdd OAI21X1
XOAI21X1_337 XOR2X1_20/Y OAI21X1_337/B OAI21X1_337/C gnd OAI21X1_337/Y vdd OAI21X1
XOAI21X1_304 AOI22X1_35/Y AOI22X1_36/Y OAI21X1_304/C gnd AOI22X1_37/D vdd OAI21X1
XNAND2X1_354 dy[12] dx[12] gnd INVX1_293/A vdd NAND2X1
XNAND2X1_332 vertices[3] cos_alpha[9] gnd XOR2X1_23/B vdd NAND2X1
XXOR2X1_26 XOR2X1_26/A XOR2X1_26/B gnd XOR2X1_26/Y vdd XOR2X1
XXOR2X1_48 XOR2X1_48/A XOR2X1_48/B gnd XOR2X1_48/Y vdd XOR2X1
XXOR2X1_37 XOR2X1_37/A XOR2X1_37/B gnd XOR2X1_37/Y vdd XOR2X1
XNAND2X1_343 AND2X2_63/Y AND2X2_76/Y gnd OAI21X1_395/C vdd NAND2X1
XNAND2X1_321 cos_gamma[3] NAND3X1_399/B gnd OR2X2_37/A vdd NAND2X1
XNAND2X1_310 INVX1_295/A NAND3X1_330/C gnd OAI21X1_363/C vdd NAND2X1
XXOR2X1_15 XOR2X1_15/A XOR2X1_15/B gnd XOR2X1_15/Y vdd XOR2X1
XNOR3X1_50 NOR3X1_50/A NOR3X1_50/B NOR3X1_50/C gnd NOR3X1_51/C vdd NOR3X1
XNAND2X1_387 vertices[4] cos_alpha[9] gnd OAI21X1_486/A vdd NAND2X1
XNAND2X1_365 OR2X2_36/B OR2X2_36/A gnd NAND2X1_366/A vdd NAND2X1
XNAND2X1_376 OAI21X1_378/Y XNOR2X1_43/Y gnd NAND3X1_436/B vdd NAND2X1
XNAND2X1_398 INVX1_316/A XOR2X1_28/Y gnd NAND3X1_408/B vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 NAND3X1_5/A NAND3X1_5/B INVX1_49/Y gnd INVX1_75/A vdd NAND3X1
XOAI21X1_112 INVX1_106/Y NOR2X1_63/A INVX1_107/A gnd XOR2X1_8/B vdd OAI21X1
XOAI21X1_101 NOR2X1_78/Y AND2X2_30/Y INVX1_127/A gnd NAND3X1_76/C vdd OAI21X1
XINVX1_209 NOR3X1_21/A gnd INVX1_209/Y vdd INVX1
XOAI21X1_178 INVX1_16/Y INVX1_146/Y OAI21X1_224/A gnd OAI21X1_179/C vdd OAI21X1
XOAI21X1_123 XNOR2X1_19/B NOR2X1_81/A INVX1_136/A gnd XNOR2X1_23/B vdd OAI21X1
XOAI21X1_134 INVX1_98/A AOI21X1_57/Y INVX1_156/A gnd OAI21X1_154/C vdd OAI21X1
XOAI21X1_156 AOI21X1_74/Y NOR3X1_15/Y INVX1_161/A gnd AOI21X1_76/A vdd OAI21X1
XOAI21X1_145 INVX1_127/A AND2X2_30/Y NAND3X1_71/C gnd AOI21X1_86/C vdd OAI21X1
XOAI21X1_189 AOI21X1_87/Y AOI21X1_88/Y OAI21X1_189/C gnd AOI21X1_91/A vdd OAI21X1
XOAI21X1_167 INVX1_168/Y XNOR2X1_30/B OAI21X1_167/C gnd NOR2X1_92/B vdd OAI21X1
XNAND2X1_173 vertices[3] cos_alpha[6] gnd OAI21X1_224/A vdd NAND2X1
XNAND2X1_151 INVX1_142/A OAI21X1_218/A gnd AOI21X1_73/A vdd NAND2X1
XNAND2X1_195 XNOR2X1_26/B XNOR2X1_26/A gnd AOI22X1_30/A vdd NAND2X1
XNAND2X1_184 INVX1_171/Y AOI22X1_31/A gnd NAND3X1_205/C vdd NAND2X1
XNAND2X1_162 OAI21X1_171/Y OR2X2_19/Y gnd OAI21X1_172/C vdd NAND2X1
XNAND2X1_140 cos_alpha[3] vertices[5] gnd OAI22X1_7/A vdd NAND2X1
XAOI22X1_18 AOI22X1_18/A AOI22X1_18/B INVX1_181/A AOI22X1_18/D gnd AOI22X1_18/Y vdd
+ AOI22X1
XAOI22X1_29 AND2X2_59/A OR2X2_25/Y INVX1_254/A AOI22X1_29/D gnd AOI22X1_29/Y vdd AOI22X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_9/C vdd NOR3X1
XXNOR2X1_84 NOR3X1_48/B INVX1_383/A gnd XNOR2X1_84/Y vdd XNOR2X1
XXNOR2X1_73 XNOR2X1_73/A XOR2X1_49/A gnd XNOR2X1_73/Y vdd XNOR2X1
XXNOR2X1_62 XNOR2X1_62/A XNOR2X1_62/B gnd INVX1_373/A vdd XNOR2X1
XXNOR2X1_51 OR2X2_56/A OR2X2_56/B gnd XOR2X1_37/A vdd XNOR2X1
XXNOR2X1_40 XNOR2X1_40/A INVX1_334/A gnd XNOR2X1_41/A vdd XNOR2X1
XAOI21X1_40 NAND3X1_49/A AOI22X1_9/D NOR3X1_4/Y gnd NOR3X1_14/C vdd AOI21X1
XAOI21X1_51 AOI21X1_51/A INVX1_93/Y NOR2X1_64/B gnd NOR3X1_10/A vdd AOI21X1
XAOI21X1_84 AOI21X1_84/A AOI21X1_84/B AOI21X1_84/C gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_95 INVX1_155/Y AOI21X1_95/B INVX1_183/Y gnd AOI21X1_95/Y vdd AOI21X1
XAOI21X1_73 AOI21X1_73/A AOI21X1_73/B INVX1_160/A gnd NOR3X1_15/C vdd AOI21X1
XAOI21X1_62 NAND3X1_76/C NAND3X1_76/A NAND3X1_72/A gnd AOI21X1_62/Y vdd AOI21X1
XOAI21X1_2 OR2X2_3/A INVX1_9/Y OAI21X1_2/C gnd NOR2X1_7/B vdd OAI21X1
XFILL_9_0_1 gnd vdd FILL
XAND2X2_109 AND2X2_109/A AND2X2_109/B gnd AND2X2_109/Y vdd AND2X2
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XNAND3X1_515 vertices[0] cos_alpha[15] INVX1_375/Y gnd NAND3X1_515/Y vdd NAND3X1
XNAND3X1_548 INVX1_386/Y NAND3X1_548/B NAND3X1_548/C gnd NAND3X1_548/Y vdd NAND3X1
XNAND3X1_537 AOI22X1_59/C AOI22X1_59/D NOR3X1_51/A gnd NAND3X1_538/C vdd NAND3X1
XNAND3X1_504 INVX1_330/Y NAND3X1_504/B OAI21X1_471/Y gnd NAND3X1_505/C vdd NAND3X1
XNAND3X1_526 INVX1_378/A NAND3X1_530/A OAI21X1_501/Y gnd NAND3X1_527/A vdd NAND3X1
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XINVX1_381 NOR3X1_48/B gnd INVX1_381/Y vdd INVX1
XFILL_24_2_2 gnd vdd FILL
XNAND3X1_345 INVX1_278/A NAND3X1_345/B OAI21X1_327/Y gnd NAND3X1_346/C vdd NAND3X1
XNAND3X1_356 NAND3X1_356/A OAI21X1_343/Y AND2X2_77/Y gnd NAND3X1_357/A vdd NAND3X1
XNAND3X1_389 INVX1_296/A NAND3X1_391/A AND2X2_94/A gnd AND2X2_95/B vdd NAND3X1
XNAND3X1_378 NAND3X1_378/A NAND3X1_378/B OAI21X1_359/Y gnd NAND3X1_379/C vdd NAND3X1
XNAND3X1_367 AND2X2_64/A OAI21X1_354/Y AND2X2_79/Y gnd NAND3X1_429/C vdd NAND3X1
XNAND3X1_312 INVX1_249/A NAND3X1_312/B NAND3X1_312/C gnd NAND3X1_315/C vdd NAND3X1
XNAND3X1_301 NAND3X1_301/A NAND3X1_301/B OAI21X1_292/C gnd NAND3X1_302/B vdd NAND3X1
XFILL_15_2_2 gnd vdd FILL
XNAND3X1_323 AOI22X1_36/C NAND3X1_323/B AOI22X1_36/D gnd NAND3X1_330/B vdd NAND3X1
XNAND3X1_334 OAI21X1_306/C NAND3X1_334/B NAND3X1_334/C gnd NAND3X1_335/B vdd NAND3X1
XOAI21X1_508 NOR3X1_49/B NOR3X1_49/C XOR2X1_52/Y gnd AOI22X1_59/D vdd OAI21X1
XNAND2X1_525 XNOR2X1_77/Y NAND2X1_525/B gnd NAND3X1_523/B vdd NAND2X1
XNAND2X1_514 XNOR2X1_67/Y NOR2X1_192/B gnd AOI22X1_57/D vdd NAND2X1
XNAND2X1_503 vertices[6] cos_alpha[9] gnd XNOR2X1_64/B vdd NAND2X1
XNAND2X1_536 cos_gamma[8] NAND2X1_536/B gnd XNOR2X1_79/B vdd NAND2X1
XAOI21X1_171 OAI21X1_395/C INVX1_288/Y INVX1_287/Y gnd NOR3X1_28/B vdd AOI21X1
XAOI21X1_182 OAI21X1_349/Y NAND3X1_362/Y INVX1_276/A gnd NOR3X1_34/C vdd AOI21X1
XAOI21X1_193 NAND3X1_396/B NAND3X1_396/C INVX1_297/A gnd AOI21X1_215/A vdd AOI21X1
XAOI21X1_160 NAND3X1_330/C NAND3X1_330/B OAI21X1_305/C gnd OAI21X1_310/B vdd AOI21X1
XNAND3X1_142 INVX1_173/A OAI21X1_153/Y AOI21X1_56/Y gnd OAI21X1_219/A vdd NAND3X1
XNAND3X1_164 AOI22X1_22/C AOI22X1_22/D AND2X2_39/Y gnd AOI21X1_75/A vdd NAND3X1
XNAND3X1_153 BUFX2_8/Y INVX1_142/A NAND3X1_457/B gnd AOI22X1_21/C vdd NAND3X1
XNAND3X1_197 INVX1_173/A INVX1_201/A OAI21X1_195/Y gnd NAND3X1_201/B vdd NAND3X1
XNAND3X1_131 AOI21X1_85/B AOI21X1_85/C AOI21X1_85/A gnd INVX1_182/A vdd NAND3X1
XNAND3X1_120 OAI21X1_177/C INVX1_150/A NAND3X1_120/C gnd NAND3X1_133/B vdd NAND3X1
XNAND3X1_186 AOI21X1_93/B AOI21X1_93/A AOI21X1_93/C gnd NAND3X1_190/C vdd NAND3X1
XNAND3X1_175 INVX1_175/A NAND3X1_184/B OAI21X1_182/Y gnd NAND3X1_175/Y vdd NAND3X1
XFILL_21_0_2 gnd vdd FILL
XOAI21X1_305 AOI22X1_35/Y AOI22X1_36/Y OAI21X1_305/C gnd OAI21X1_305/Y vdd OAI21X1
XOAI21X1_327 INVX1_45/Y INVX1_241/Y XOR2X1_23/Y gnd OAI21X1_327/Y vdd OAI21X1
XOAI21X1_349 NOR3X1_35/B NOR3X1_35/C OAI21X1_349/C gnd OAI21X1_349/Y vdd OAI21X1
XOAI21X1_338 INVX1_286/A AND2X2_75/Y INVX1_285/Y gnd AND2X2_77/B vdd OAI21X1
XOAI21X1_316 INVX1_229/Y NOR2X1_133/A OAI21X1_316/C gnd AND2X2_71/B vdd OAI21X1
XXOR2X1_27 OR2X2_38/A OR2X2_38/B gnd XOR2X1_27/Y vdd XOR2X1
XNAND2X1_333 NOR2X1_141/Y XOR2X1_23/Y gnd NAND3X1_344/C vdd NAND2X1
XXOR2X1_38 OR2X2_53/A OR2X2_53/B gnd XOR2X1_38/Y vdd XOR2X1
XXOR2X1_49 XOR2X1_49/A XOR2X1_49/B gnd XOR2X1_49/Y vdd XOR2X1
XNAND2X1_377 AND2X2_89/Y XOR2X1_26/Y gnd NAND3X1_436/C vdd NAND2X1
XNAND2X1_300 dy[11] dx[11] gnd INVX1_251/A vdd NAND2X1
XNAND2X1_366 NAND2X1_366/A OR2X2_36/Y gnd INVX1_306/A vdd NAND2X1
XNAND2X1_355 AND2X2_87/A NAND3X1_376/Y gnd NAND3X1_379/A vdd NAND2X1
XNAND2X1_344 BUFX2_16/Y vertices[12] gnd OR2X2_40/A vdd NAND2X1
XNAND2X1_322 OR2X2_37/B OR2X2_37/A gnd OAI21X1_321/C vdd NAND2X1
XNAND2X1_311 cos_gamma[6] NOR2X1_73/Y gnd NOR2X1_166/A vdd NAND2X1
XXOR2X1_16 XOR2X1_16/A XOR2X1_16/B gnd XOR2X1_16/Y vdd XOR2X1
XNOR3X1_51 NOR3X1_51/A NOR3X1_51/B NOR3X1_51/C gnd NOR3X1_51/Y vdd NOR3X1
XNOR3X1_40 NOR3X1_40/A NOR3X1_40/B NOR3X1_40/C gnd NOR3X1_41/C vdd NOR3X1
XNAND2X1_388 vertices[4] cos_alpha[10] gnd OAI21X1_437/C vdd NAND2X1
XNAND2X1_399 OAI21X1_394/Y OR2X2_39/Y gnd OAI21X1_440/A vdd NAND2X1
XFILL_4_1_2 gnd vdd FILL
XFILL_12_0_2 gnd vdd FILL
XNAND3X1_6 INVX1_47/Y INVX1_75/A NAND3X1_6/C gnd INVX1_53/A vdd NAND3X1
XOAI21X1_113 NOR3X1_5/B NOR3X1_5/C NOR3X1_5/A gnd AOI21X1_48/A vdd OAI21X1
XOAI21X1_135 NAND3X1_80/A AOI21X1_58/Y NAND3X1_82/B gnd AOI21X1_84/C vdd OAI21X1
XOAI21X1_124 INVX1_92/Y NOR3X1_11/B AOI21X1_53/B gnd INVX1_137/A vdd OAI21X1
XOAI21X1_102 INVX1_1/Y INVX1_128/Y NOR2X1_78/A gnd NAND3X1_71/B vdd OAI21X1
XOAI21X1_146 INVX1_1/Y OAI22X1_6/D OAI21X1_146/C gnd AOI22X1_24/D vdd OAI21X1
XOAI21X1_157 NOR3X1_15/B NOR3X1_15/C NOR3X1_15/A gnd OAI21X1_157/Y vdd OAI21X1
XOAI21X1_168 NOR2X1_91/A NOR2X1_7/B NOR2X1_92/B gnd OAI21X1_168/Y vdd OAI21X1
XOAI21X1_179 INVX1_147/A INVX1_205/A OAI21X1_179/C gnd OR2X2_22/A vdd OAI21X1
XNAND2X1_152 dy[8] dx[8] gnd INVX1_158/A vdd NAND2X1
XNAND2X1_130 OAI21X1_169/A AND2X2_36/Y gnd NAND3X1_114/C vdd NAND2X1
XNAND2X1_185 NAND3X1_202/C NAND2X1_185/B gnd NAND3X1_204/C vdd NAND2X1
XNAND2X1_163 OR2X2_20/B OR2X2_20/A gnd OAI21X1_213/C vdd NAND2X1
XNAND2X1_196 AND2X2_56/B AND2X2_56/A gnd OAI21X1_250/C vdd NAND2X1
XNAND2X1_141 AOI22X1_18/A AOI22X1_18/B gnd AOI21X1_66/C vdd NAND2X1
XNAND2X1_174 vertices[1] cos_alpha[8] gnd OR2X2_22/B vdd NAND2X1
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XAOI22X1_19 AOI22X1_19/A AOI22X1_19/B INVX1_182/A AOI22X1_19/D gnd AOI22X1_19/Y vdd
+ AOI22X1
XXNOR2X1_41 XNOR2X1_41/A XNOR2X1_41/B gnd OR2X2_36/A vdd XNOR2X1
XXNOR2X1_30 INVX1_229/A XNOR2X1_30/B gnd INVX1_197/A vdd XNOR2X1
XXNOR2X1_63 XNOR2X1_63/A XNOR2X1_63/B gnd XNOR2X1_63/Y vdd XNOR2X1
XXNOR2X1_74 XOR2X1_48/Y XOR2X1_49/A gnd XNOR2X1_74/Y vdd XNOR2X1
XXNOR2X1_52 XOR2X1_37/Y XNOR2X1_52/B gnd OR2X2_53/A vdd XNOR2X1
XAOI21X1_52 AOI21X1_52/A AOI21X1_52/B INVX1_133/Y gnd NOR3X1_10/B vdd AOI21X1
XAOI21X1_30 NAND2X1_99/B OAI21X1_84/Y INVX1_90/A gnd NOR3X1_12/B vdd AOI21X1
XAOI21X1_41 NOR2X1_59/Y OAI21X1_77/Y NOR3X1_3/Y gnd NAND3X1_85/C vdd AOI21X1
XOAI21X1_3 INVX1_3/A INVX1_11/Y OAI22X1_1/Y gnd OAI21X1_5/A vdd OAI21X1
XAOI21X1_74 AOI21X1_74/A AOI21X1_74/B XOR2X1_10/Y gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_85 AOI21X1_85/A AOI21X1_85/B AOI21X1_85/C gnd AOI21X1_85/Y vdd AOI21X1
XFILL_9_0_2 gnd vdd FILL
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B AND2X2_45/Y gnd AOI21X1_96/Y vdd AOI21X1
XAOI21X1_63 AOI21X1_63/A AOI21X1_63/B INVX1_154/A gnd AOI21X1_63/Y vdd AOI21X1
XFILL_27_2_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A XOR2X1_6/B gnd XOR2X1_6/Y vdd XOR2X1
XNAND3X1_538 INVX1_380/Y INVX1_381/Y NAND3X1_538/C gnd NAND3X1_539/B vdd NAND3X1
XNAND3X1_516 INVX1_376/A OAI21X1_490/Y NAND3X1_516/C gnd NAND3X1_519/B vdd NAND3X1
XNAND3X1_505 NAND3X1_505/A NAND3X1_505/B NAND3X1_505/C gnd AOI22X1_56/B vdd NAND3X1
XNAND3X1_527 NAND3X1_527/A OAI21X1_502/Y NOR3X1_46/Y gnd NAND3X1_532/A vdd NAND3X1
XFILL_10_1_0 gnd vdd FILL
XFILL_18_2_0 gnd vdd FILL
XINVX1_360 dz[14] gnd INVX1_360/Y vdd INVX1
XINVX1_382 NOR3X1_50/B gnd INVX1_382/Y vdd INVX1
XINVX1_371 XOR2X1_34/B gnd INVX1_371/Y vdd INVX1
XNAND3X1_346 INVX1_309/A NAND3X1_346/B NAND3X1_346/C gnd INVX1_280/A vdd NAND3X1
XNAND3X1_357 NAND3X1_357/A OAI21X1_337/Y OAI21X1_342/Y gnd OAI21X1_389/C vdd NAND3X1
XNAND3X1_379 NAND3X1_379/A NAND3X1_379/B NAND3X1_379/C gnd NAND3X1_383/A vdd NAND3X1
XNAND3X1_368 INVX1_273/Y NAND3X1_368/B OAI21X1_355/Y gnd NAND3X1_373/C vdd NAND3X1
XNAND3X1_313 BUFX2_7/Y AOI22X1_31/B AOI22X1_45/B gnd NAND3X1_314/B vdd NAND3X1
XNAND3X1_302 INVX1_240/A NAND3X1_302/B OAI21X1_293/Y gnd NAND3X1_306/C vdd NAND3X1
XNAND3X1_324 INVX1_234/Y AND2X2_67/B NAND3X1_324/C gnd AOI22X1_36/A vdd NAND3X1
XNAND3X1_335 INVX1_256/Y NAND3X1_335/B OAI21X1_307/Y gnd AOI22X1_39/D vdd NAND3X1
XOAI21X1_509 OAI21X1_509/A NOR3X1_48/Y INVX1_368/Y gnd AOI22X1_60/D vdd OAI21X1
XFILL_15_1 gnd vdd FILL
XNAND2X1_526 NAND3X1_521/Y NAND3X1_523/Y gnd NAND3X1_524/C vdd NAND2X1
XNAND2X1_504 vertices[4] cos_alpha[11] gnd XNOR2X1_65/B vdd NAND2X1
XNAND2X1_515 XOR2X1_49/B XNOR2X1_74/Y gnd AOI22X1_57/A vdd NAND2X1
XNAND2X1_537 OR2X2_59/B OR2X2_59/A gnd NAND3X1_534/A vdd NAND2X1
XINVX1_190 INVX1_190/A gnd INVX1_190/Y vdd INVX1
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 INVX1_202/Y OAI21X1_239/Y INVX1_248/Y gnd OAI21X1_295/C vdd AOI21X1
XAOI21X1_183 NAND3X1_362/C OAI21X1_347/Y OAI21X1_349/C gnd OAI21X1_379/B vdd AOI21X1
XAOI21X1_172 OAI21X1_341/Y NAND3X1_412/B OAI21X1_340/Y gnd NOR3X1_29/A vdd AOI21X1
XAOI21X1_194 NOR2X1_152/B NOR2X1_152/A AOI21X1_215/A gnd XOR2X1_32/B vdd AOI21X1
XAOI21X1_161 AOI22X1_33/D NAND3X1_321/B INVX1_270/Y gnd INVX1_271/A vdd AOI21X1
XFILL_7_1_0 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XNAND3X1_110 OAI21X1_87/Y AOI21X1_54/B AOI21X1_54/A gnd AOI21X1_53/B vdd NAND3X1
XNAND3X1_121 INVX1_151/Y NAND3X1_133/B OAI21X1_140/Y gnd AOI22X1_19/B vdd NAND3X1
XNAND3X1_132 INVX1_151/Y NAND3X1_132/B OAI21X1_139/Y gnd AOI22X1_20/A vdd NAND3X1
XNAND3X1_143 NAND3X1_96/C INVX1_173/A OAI21X1_153/Y gnd NAND3X1_151/B vdd NAND3X1
XNAND3X1_165 INVX1_163/A AOI21X1_75/B AOI21X1_75/A gnd INVX1_162/A vdd NAND3X1
XNAND3X1_154 OAI21X1_219/A AOI21X1_72/Y NAND3X1_154/C gnd NOR2X1_107/A vdd NAND3X1
XNAND3X1_198 NAND3X1_198/A OAI21X1_196/Y INVX1_173/Y gnd NAND3X1_201/C vdd NAND3X1
XNAND3X1_187 INVX1_213/A AOI21X1_92/A AOI21X1_92/C gnd NAND3X1_190/A vdd NAND3X1
XNAND3X1_176 INVX1_178/A AOI21X1_88/A AOI21X1_88/B gnd NAND3X1_180/A vdd NAND3X1
XOAI21X1_328 NOR2X1_121/Y INVX1_281/Y OAI21X1_328/C gnd OAI21X1_329/C vdd OAI21X1
XOAI21X1_317 NOR2X1_83/A OAI22X1_8/D NOR2X1_166/A gnd INVX1_266/A vdd OAI21X1
XOAI21X1_306 AOI22X1_37/Y OAI21X1_307/B OAI21X1_306/C gnd AOI22X1_38/D vdd OAI21X1
XOAI21X1_339 INVX1_28/Y OAI22X1_6/B AND2X2_75/A gnd OAI21X1_339/Y vdd OAI21X1
XNAND2X1_389 INVX1_312/Y XOR2X1_27/Y gnd NAND3X1_402/B vdd NAND2X1
XXOR2X1_39 XOR2X1_39/A XOR2X1_39/B gnd XOR2X1_39/Y vdd XOR2X1
XNAND2X1_334 vertices[3] cos_alpha[10] gnd OAI21X1_325/B vdd NAND2X1
XXOR2X1_17 XOR2X1_17/A XOR2X1_17/B gnd XOR2X1_17/Y vdd XOR2X1
XNAND2X1_367 INVX1_303/Y XNOR2X1_42/Y gnd AOI22X1_48/A vdd NAND2X1
XNAND2X1_378 XNOR2X1_43/Y AND2X2_89/Y gnd NAND3X1_437/C vdd NAND2X1
XNAND2X1_345 AND2X2_74/B AND2X2_74/A gnd NOR3X1_31/B vdd NAND2X1
XXOR2X1_28 OR2X2_39/A OR2X2_39/B gnd XOR2X1_28/Y vdd XOR2X1
XNAND2X1_356 AOI22X1_44/A AOI22X1_44/B gnd NOR2X1_152/A vdd NAND2X1
XNAND2X1_312 OR2X2_30/B OR2X2_30/A gnd AND2X2_70/B vdd NAND2X1
XNAND2X1_323 cos_gamma[4] NAND3X1_399/B gnd OAI21X1_377/C vdd NAND2X1
XNAND2X1_301 AND2X2_72/A AOI22X1_33/B gnd NAND3X1_320/B vdd NAND2X1
XNOR3X1_52 NOR3X1_52/A NOR3X1_52/B NOR3X1_52/C gnd NOR3X1_52/Y vdd NOR3X1
XNOR3X1_41 NOR3X1_41/A NOR3X1_41/B NOR3X1_41/C gnd NOR3X1_41/Y vdd NOR3X1
XNOR3X1_30 NOR3X1_30/A NOR3X1_30/B NOR3X1_30/C gnd NOR3X1_31/C vdd NOR3X1
XNAND3X1_7 NOR3X1_2/B INVX1_53/A INVX1_54/Y gnd NAND3X1_8/B vdd NAND3X1
XOAI21X1_114 NOR3X1_6/B NOR3X1_6/C NOR3X1_6/A gnd AOI21X1_47/A vdd OAI21X1
XOAI21X1_125 NOR3X1_9/A NOR3X1_9/B AOI21X1_52/B gnd INVX1_164/A vdd OAI21X1
XOAI21X1_103 NOR3X1_13/A NOR3X1_13/B NOR3X1_13/C gnd NAND3X1_78/C vdd OAI21X1
XOAI21X1_158 AOI21X1_74/Y NOR3X1_15/Y INVX1_161/Y gnd AOI22X1_22/D vdd OAI21X1
XOAI21X1_169 OAI21X1_169/A AND2X2_36/Y AND2X2_39/A gnd XNOR2X1_26/A vdd OAI21X1
XOAI21X1_147 AOI21X1_63/Y AOI22X1_17/Y AOI21X1_86/C gnd AOI21X1_66/A vdd OAI21X1
XOAI21X1_136 INVX1_45/Y INVX1_146/Y INVX1_147/Y gnd AOI21X1_61/A vdd OAI21X1
XBUFX2_1 cos_alpha[0] gnd INVX1_1/A vdd BUFX2
XNAND2X1_164 XOR2X1_10/B XOR2X1_10/A gnd NAND2X1_165/A vdd NAND2X1
XNAND2X1_197 INVX1_193/Y XNOR2X1_25/A gnd NAND2X1_198/B vdd NAND2X1
XNAND2X1_120 NAND3X1_75/Y AOI22X1_13/B gnd NAND3X1_78/B vdd NAND2X1
XNAND2X1_153 AOI21X1_81/A INVX1_166/Y gnd XNOR2X1_23/A vdd NAND2X1
XNAND2X1_131 AND2X2_35/Y AND2X2_36/Y gnd NAND3X1_115/C vdd NAND2X1
XNAND2X1_186 INVX1_171/A NAND3X1_204/Y gnd NAND3X1_205/B vdd NAND2X1
XNAND2X1_175 NAND3X1_173/Y NAND3X1_175/Y gnd AOI21X1_92/C vdd NAND2X1
XNAND2X1_142 NOR2X1_97/A NOR2X1_97/B gnd AOI22X1_17/D vdd NAND2X1
XAOI21X1_1 XOR2X1_4/B AOI21X1_1/B INVX1_34/Y gnd INVX1_35/A vdd AOI21X1
XXNOR2X1_53 XNOR2X1_53/A INVX1_360/Y gnd XOR2X1_39/A vdd XNOR2X1
XXNOR2X1_64 XNOR2X1_64/A XNOR2X1_64/B gnd XNOR2X1_65/A vdd XNOR2X1
XXNOR2X1_75 XOR2X1_49/A XOR2X1_49/B gnd XNOR2X1_75/Y vdd XNOR2X1
XXNOR2X1_42 XNOR2X1_42/A INVX1_306/A gnd XNOR2X1_42/Y vdd XNOR2X1
XXNOR2X1_20 XOR2X1_9/Y NOR2X1_82/Y gnd NOR2X1_84/A vdd XNOR2X1
XXNOR2X1_31 XNOR2X1_31/A XNOR2X1_31/B gnd OR2X2_25/A vdd XNOR2X1
XBUFX2_30 BUFX2_30/A gnd vertices_out[12] vdd BUFX2
XAOI21X1_42 NAND3X1_80/C NAND3X1_80/B NAND3X1_80/A gnd AOI21X1_42/Y vdd AOI21X1
XAOI21X1_53 AOI21X1_53/A AOI21X1_53/B INVX1_92/A gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_20 OAI21X1_47/Y INVX1_76/A OAI21X1_51/C gnd OAI21X1_67/B vdd AOI21X1
XAOI21X1_31 INVX1_94/A NAND3X1_34/B NOR2X1_55/Y gnd NOR2X1_69/B vdd AOI21X1
XAOI21X1_75 AOI21X1_75/A AOI21X1_75/B INVX1_163/A gnd AOI21X1_75/Y vdd AOI21X1
XAOI21X1_64 NAND3X1_71/B INVX1_127/Y NOR2X1_78/Y gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_86 AOI21X1_86/A AOI21X1_86/B AOI21X1_86/C gnd AOI21X1_86/Y vdd AOI21X1
XOAI21X1_4 INVX1_4/Y INVX1_5/Y AND2X2_1/B gnd XNOR2X1_1/B vdd OAI21X1
XAOI21X1_97 AOI21X1_97/A AOI21X1_97/B AOI21X1_97/C gnd AOI21X1_97/Y vdd AOI21X1
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A XOR2X1_7/B gnd XOR2X1_7/Y vdd XOR2X1
XNAND3X1_539 INVX1_368/A NAND3X1_539/B OAI21X1_510/Y gnd AOI22X1_60/C vdd NAND3X1
XNAND3X1_517 NAND3X1_517/A OAI21X1_493/Y OAI21X1_494/Y gnd NAND3X1_518/B vdd NAND3X1
XNAND3X1_506 AOI22X1_54/C NAND3X1_506/B AOI22X1_54/D gnd OAI21X1_479/C vdd NAND3X1
XNAND3X1_528 INVX1_377/A NAND3X1_528/B AND2X2_108/Y gnd NAND3X1_529/C vdd NAND3X1
XFILL_10_1_1 gnd vdd FILL
XFILL_18_2_1 gnd vdd FILL
XINVX1_383 INVX1_383/A gnd INVX1_383/Y vdd INVX1
XINVX1_361 INVX1_361/A gnd INVX1_361/Y vdd INVX1
XINVX1_350 cos_alpha[14] gnd INVX1_350/Y vdd INVX1
XINVX1_372 XOR2X1_49/B gnd INVX1_372/Y vdd INVX1
XNAND3X1_314 INVX1_249/Y NAND3X1_314/B NAND3X1_314/C gnd NAND3X1_315/B vdd NAND3X1
XNAND3X1_303 INVX1_240/Y INVX1_274/A OAI21X1_292/Y gnd NAND3X1_306/B vdd NAND3X1
XNAND3X1_347 INVX1_280/A OAI21X1_330/C INVX1_279/Y gnd NAND3X1_348/C vdd NAND3X1
XNAND3X1_358 OAI21X1_389/C OAI21X1_344/Y AND2X2_74/Y gnd NAND3X1_359/B vdd NAND3X1
XNAND3X1_369 BUFX2_9/Y OAI21X1_355/C NAND3X1_369/C gnd AND2X2_89/B vdd NAND3X1
XNAND3X1_325 INVX1_234/A NAND3X1_325/B NAND3X1_325/C gnd AOI22X1_36/B vdd NAND3X1
XNAND3X1_336 INVX1_256/Y INVX1_297/A AOI22X1_38/D gnd OAI21X1_366/C vdd NAND3X1
XFILL_15_2 gnd vdd FILL
XNAND2X1_527 INVX1_349/Y XNOR2X1_48/A gnd OR2X2_58/B vdd NAND2X1
XNAND2X1_516 INVX1_372/Y XNOR2X1_73/Y gnd AOI22X1_57/B vdd NAND2X1
XNAND2X1_505 XOR2X1_36/B XOR2X1_36/A gnd AND2X2_105/A vdd NAND2X1
XNAND2X1_538 NAND3X1_534/A OR2X2_59/Y gnd NAND2X1_539/B vdd NAND2X1
XINVX1_191 INVX1_191/A gnd NOR3X1_22/B vdd INVX1
XINVX1_180 OAI22X1_7/C gnd INVX1_180/Y vdd INVX1
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_184 OAI21X1_350/Y NAND3X1_364/A INVX1_290/Y gnd OAI21X1_351/A vdd AOI21X1
XAOI21X1_140 OAI21X1_284/Y OAI21X1_337/C XNOR2X1_34/Y gnd NOR3X1_24/B vdd AOI21X1
XAOI21X1_173 XNOR2X1_34/Y OAI21X1_284/Y NOR3X1_23/Y gnd NOR3X1_30/B vdd AOI21X1
XAOI21X1_162 INVX1_249/Y NAND3X1_314/C NOR2X1_137/Y gnd OAI21X1_375/B vdd AOI21X1
XAOI21X1_151 NAND3X1_252/C NAND3X1_252/B INVX1_201/A gnd NAND3X1_307/A vdd AOI21X1
XAOI21X1_195 NOR2X1_136/Y INVX1_267/A AND2X2_71/Y gnd INVX1_303/A vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XNAND3X1_111 INVX1_92/A AOI21X1_53/B AOI21X1_53/A gnd NAND3X1_112/A vdd NAND3X1
XNAND3X1_100 NAND3X1_95/A NAND3X1_98/B NAND3X1_98/C gnd NAND3X1_101/C vdd NAND3X1
XNAND3X1_144 NAND3X1_144/A NAND3X1_144/B AOI21X1_68/Y gnd AOI21X1_83/B vdd NAND3X1
XNAND3X1_166 INVX1_140/A INVX1_162/A AOI21X1_77/A gnd INVX1_165/A vdd NAND3X1
XNAND3X1_155 NAND3X1_99/Y NAND3X1_155/B NAND3X1_155/C gnd NAND3X1_156/C vdd NAND3X1
XNAND3X1_133 NOR2X1_75/B NAND3X1_133/B OAI21X1_140/Y gnd AOI22X1_20/B vdd NAND3X1
XNAND3X1_122 NOR2X1_87/Y AOI22X1_23/D NAND3X1_122/C gnd AOI22X1_18/A vdd NAND3X1
XNAND3X1_177 INVX1_178/Y OAI22X1_6/Y AOI21X1_87/A gnd NAND3X1_180/B vdd NAND3X1
XNAND3X1_199 NAND3X1_200/A NAND3X1_201/B NAND3X1_201/C gnd NAND3X1_199/Y vdd NAND3X1
XNAND3X1_188 NAND3X1_190/A NAND3X1_190/C AOI21X1_94/Y gnd AOI21X1_97/A vdd NAND3X1
XOAI21X1_329 INVX1_279/A INVX1_280/Y OAI21X1_329/C gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_318 NOR2X1_136/A AND2X2_71/Y INVX1_267/Y gnd OAI21X1_318/Y vdd OAI21X1
XOAI21X1_307 AOI22X1_37/Y OAI21X1_307/B OAI21X1_307/C gnd OAI21X1_307/Y vdd OAI21X1
XXOR2X1_18 XOR2X1_18/A XOR2X1_18/B gnd XOR2X1_18/Y vdd XOR2X1
XNAND2X1_302 AOI22X1_34/A AOI22X1_34/B gnd NAND3X1_321/B vdd NAND2X1
XNAND2X1_335 NOR2X1_141/Y OAI21X1_326/C gnd NAND3X1_345/B vdd NAND2X1
XNAND2X1_357 AND2X2_95/B AND2X2_95/A gnd NAND3X1_453/A vdd NAND2X1
XNOR3X1_42 NOR3X1_42/A NOR3X1_42/B NOR3X1_42/C gnd NOR3X1_42/Y vdd NOR3X1
XNOR3X1_31 NOR3X1_31/A NOR3X1_31/B NOR3X1_31/C gnd NOR3X1_32/C vdd NOR3X1
XXOR2X1_29 XOR2X1_29/A OR2X2_57/A gnd XOR2X1_30/A vdd XOR2X1
XNAND2X1_368 INVX1_306/Y XNOR2X1_42/A gnd OAI21X1_418/C vdd NAND2X1
XNAND2X1_379 OAI21X1_378/Y XOR2X1_26/Y gnd NAND3X1_437/B vdd NAND2X1
XNAND2X1_313 INVX1_267/A NOR2X1_136/Y gnd NAND2X1_314/B vdd NAND2X1
XNAND2X1_346 INVX1_359/A AND2X2_79/A gnd OAI21X1_406/A vdd NAND2X1
XNAND2X1_324 OAI21X1_375/B XNOR2X1_38/Y gnd NAND3X1_375/B vdd NAND2X1
XNOR3X1_20 NOR3X1_20/A NOR3X1_20/B NOR3X1_20/C gnd NOR3X1_20/Y vdd NOR3X1
XNAND3X1_8 NAND3X1_8/A NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_115 INVX1_110/Y NAND2X1_97/B INVX1_118/A gnd AOI21X1_49/C vdd OAI21X1
XOAI21X1_104 NOR2X1_76/Y NOR2X1_77/Y INVX1_126/Y gnd AOI22X1_13/B vdd OAI21X1
XOAI21X1_159 AOI21X1_75/Y INVX1_162/Y INVX1_140/Y gnd AOI21X1_79/A vdd OAI21X1
XOAI21X1_148 AOI21X1_63/Y AOI22X1_17/Y AOI21X1_64/Y gnd AOI22X1_18/D vdd OAI21X1
XOAI21X1_126 INVX1_91/Y INVX1_18/Y NOR2X1_82/B gnd OAI21X1_127/C vdd OAI21X1
XOAI21X1_137 INVX1_16/Y INVX1_148/Y INVX1_149/Y gnd AOI21X1_61/B vdd OAI21X1
XNAND2X1_110 OR2X2_15/B OR2X2_15/A gnd INVX1_155/A vdd NAND2X1
XNAND2X1_121 INVX1_129/Y INVX1_142/A gnd AND2X2_36/B vdd NAND2X1
XNAND2X1_132 OAI21X1_169/A OAI21X1_133/Y gnd NAND3X1_115/B vdd NAND2X1
XBUFX2_2 cos_alpha[0] gnd BUFX2_2/Y vdd BUFX2
XNAND2X1_143 BUFX2_16/Y vertices[7] gnd OAI21X1_146/C vdd NAND2X1
XNAND2X1_165 NAND2X1_165/A NAND3X1_163/B gnd INVX1_188/A vdd NAND2X1
XNAND2X1_154 NOR2X1_82/Y XOR2X1_9/Y gnd OR2X2_17/B vdd NAND2X1
XNAND2X1_187 AOI21X1_98/B AOI21X1_98/A gnd NAND3X1_399/B vdd NAND2X1
XNAND2X1_176 vertices[4] cos_alpha[5] gnd OAI22X1_7/C vdd NAND2X1
XNAND2X1_198 NAND3X1_221/Y NAND2X1_198/B gnd OR2X2_25/B vdd NAND2X1
XAOI21X1_2 INVX1_30/A AOI21X1_2/B NOR2X1_25/A gnd NOR3X1_2/B vdd AOI21X1
XXNOR2X1_76 XOR2X1_44/A XOR2X1_44/B gnd XNOR2X1_76/Y vdd XNOR2X1
XXNOR2X1_65 XNOR2X1_65/A XNOR2X1_65/B gnd XNOR2X1_66/B vdd XNOR2X1
XXNOR2X1_43 XOR2X1_26/A XOR2X1_26/B gnd XNOR2X1_43/Y vdd XNOR2X1
XXNOR2X1_54 XNOR2X1_54/A XOR2X1_40/Y gnd XOR2X1_41/A vdd XNOR2X1
XXNOR2X1_32 XOR2X1_14/A XOR2X1_14/B gnd XNOR2X1_32/Y vdd XNOR2X1
XXNOR2X1_10 XNOR2X1_9/Y INVX1_21/Y gnd XNOR2X1_10/Y vdd XNOR2X1
XXNOR2X1_21 XNOR2X1_21/A NOR2X1_87/Y gnd XNOR2X1_21/Y vdd XNOR2X1
XBUFX2_31 BUFX2_31/A gnd vertices_out[13] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd vertices_out[2] vdd BUFX2
XAOI21X1_54 AOI21X1_54/A AOI21X1_54/B OAI21X1_87/Y gnd NOR3X1_11/B vdd AOI21X1
XAOI21X1_32 INVX1_110/A OAI21X1_83/Y INVX1_118/Y gnd NOR3X1_8/B vdd AOI21X1
XOAI21X1_5 OAI21X1_5/A XNOR2X1_1/Y OAI21X1_5/C gnd XOR2X1_2/B vdd OAI21X1
XAOI21X1_21 NAND3X1_20/B OAI21X1_49/Y NOR3X1_1/Y gnd NOR3X1_3/C vdd AOI21X1
XAOI21X1_65 NAND3X1_78/B NAND3X1_78/C NOR3X1_13/Y gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_10 NAND3X1_5/B NAND3X1_5/A INVX1_49/Y gnd OAI21X1_40/B vdd AOI21X1
XAOI21X1_43 NAND3X1_95/Y NAND3X1_98/Y INVX1_7/Y gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_76 AOI21X1_76/A AOI21X1_76/B AOI21X1_76/C gnd AOI21X1_76/Y vdd AOI21X1
XAOI21X1_98 AOI21X1_98/A AOI21X1_98/B INVX1_7/Y gnd AOI22X1_31/A vdd AOI21X1
XAOI21X1_87 AOI21X1_87/A OAI22X1_6/Y INVX1_178/Y gnd AOI21X1_87/Y vdd AOI21X1
XOAI21X1_490 AOI22X1_58/Y AOI22X1_57/Y INVX1_373/Y gnd OAI21X1_490/Y vdd OAI21X1
XFILL_27_2_2 gnd vdd FILL
XFILL_2_2_2 gnd vdd FILL
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B gnd XOR2X1_8/Y vdd XOR2X1
XNAND3X1_518 INVX1_376/Y NAND3X1_518/B OAI22X1_12/Y gnd NAND3X1_519/A vdd NAND3X1
XNAND3X1_507 cos_gamma[1] NAND3X1_507/B NAND3X1_528/B gnd OAI21X1_480/B vdd NAND3X1
XNAND3X1_529 INVX1_7/A OAI21X1_503/Y NAND3X1_529/C gnd NAND3X1_531/A vdd NAND3X1
XFILL_10_1_2 gnd vdd FILL
XFILL_18_2_2 gnd vdd FILL
XINVX1_351 INVX1_351/A gnd INVX1_351/Y vdd INVX1
XINVX1_384 NOR3X1_52/A gnd INVX1_384/Y vdd INVX1
XINVX1_373 INVX1_373/A gnd INVX1_373/Y vdd INVX1
XINVX1_362 XOR2X1_39/Y gnd INVX1_362/Y vdd INVX1
XINVX1_340 INVX1_340/A gnd INVX1_340/Y vdd INVX1
XDFFPOSX1_10 BUFX2_27/A clk XOR2X1_12/Y gnd vdd DFFPOSX1
XNAND3X1_337 XNOR2X1_23/B AOI22X1_39/Y NOR2X1_129/Y gnd AOI22X1_44/C vdd NAND3X1
XNAND3X1_348 INVX1_242/Y OAI21X1_329/Y NAND3X1_348/C gnd NAND3X1_348/Y vdd NAND3X1
XNAND3X1_315 XOR2X1_21/Y NAND3X1_315/B NAND3X1_315/C gnd AND2X2_80/A vdd NAND3X1
XNAND3X1_304 NAND3X1_306/C NAND3X1_306/B OAI21X1_295/C gnd NAND3X1_305/B vdd NAND3X1
XNAND3X1_326 NAND3X1_326/A NAND3X1_326/B OAI21X1_302/C gnd INVX1_295/A vdd NAND3X1
XNAND3X1_359 OAI21X1_331/Y NAND3X1_359/B OAI21X1_345/Y gnd OAI21X1_380/C vdd NAND3X1
XINVX1_170 NOR2X1_92/Y gnd INVX1_170/Y vdd INVX1
XNAND2X1_528 OR2X2_58/B OR2X2_58/A gnd NAND3X1_524/A vdd NAND2X1
XNAND2X1_517 XOR2X1_45/Y NOR2X1_192/B gnd AOI22X1_58/C vdd NAND2X1
XNAND2X1_506 AND2X2_105/B AND2X2_105/A gnd NOR2X1_191/A vdd NAND2X1
XNAND2X1_539 INVX1_379/Y NAND2X1_539/B gnd AND2X2_109/A vdd NAND2X1
XINVX1_192 INVX1_192/A gnd NOR3X1_22/C vdd INVX1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XFILL_24_0_2 gnd vdd FILL
XAOI21X1_174 OAI21X1_343/Y NAND3X1_356/A AND2X2_77/Y gnd NOR3X1_30/A vdd AOI21X1
XAOI21X1_196 NAND3X1_308/Y OAI21X1_296/Y INVX1_41/Y gnd INVX1_308/A vdd AOI21X1
XAOI21X1_185 NAND3X1_308/Y OAI21X1_296/Y INVX1_8/Y gnd OAI21X1_355/C vdd AOI21X1
XAOI21X1_141 OAI21X1_331/C OAI21X1_287/Y NAND3X1_295/C gnd OAI21X1_291/B vdd AOI21X1
XAOI21X1_163 INVX1_240/Y OAI21X1_292/Y INVX1_274/Y gnd NOR3X1_34/A vdd AOI21X1
XAOI21X1_152 NAND3X1_314/C NAND3X1_314/B INVX1_249/Y gnd NOR3X1_25/B vdd AOI21X1
XAOI21X1_130 NAND3X1_244/B NAND3X1_244/A INVX1_215/A gnd OAI21X1_266/B vdd AOI21X1
XFILL_7_1_2 gnd vdd FILL
XFILL_15_0_2 gnd vdd FILL
XNAND3X1_112 NAND3X1_112/A NOR3X1_12/C OAI21X1_122/Y gnd NOR3X1_19/A vdd NAND3X1
XNAND3X1_145 AOI21X1_71/Y AOI21X1_83/B AOI21X1_83/A gnd NAND3X1_151/C vdd NAND3X1
XNAND3X1_101 BUFX2_7/Y NAND3X1_99/Y NAND3X1_101/C gnd OAI21X1_173/A vdd NAND3X1
XNAND3X1_167 INVX1_164/A INVX1_165/A AOI21X1_79/A gnd AOI21X1_78/B vdd NAND3X1
XNAND3X1_156 BUFX2_9/Y NOR2X1_107/A NAND3X1_156/C gnd OAI21X1_218/A vdd NAND3X1
XNAND3X1_134 AOI21X1_85/B AOI21X1_85/A AOI21X1_65/Y gnd AOI22X1_20/D vdd NAND3X1
XNAND3X1_189 AOI21X1_97/C AOI21X1_97/B AOI21X1_97/A gnd NAND3X1_194/A vdd NAND3X1
XNAND3X1_123 BUFX2_3/Y vertices[8] OAI21X1_146/C gnd AOI21X1_63/A vdd NAND3X1
XNAND3X1_178 AOI22X1_24/Y NAND3X1_180/B NAND3X1_180/A gnd AOI21X1_91/B vdd NAND3X1
XFILL_20_1 gnd vdd FILL
XOAI21X1_308 INVX1_166/Y OAI21X1_308/B OAI21X1_308/C gnd OAI21X1_308/Y vdd OAI21X1
XOAI21X1_319 INVX1_236/A INVX1_237/A AND2X2_72/A gnd OAI21X1_319/Y vdd OAI21X1
XNAND2X1_336 NAND3X1_348/Y NAND3X1_350/Y gnd NOR3X1_33/A vdd NAND2X1
XXOR2X1_19 XOR2X1_19/A XOR2X1_19/B gnd XOR2X1_19/Y vdd XOR2X1
XNAND2X1_314 OAI21X1_318/Y NAND2X1_314/B gnd INVX1_268/A vdd NAND2X1
XNAND2X1_325 OAI21X1_375/B XOR2X1_22/Y gnd NAND3X1_376/B vdd NAND2X1
XNAND2X1_303 AOI22X1_36/A AOI22X1_36/B gnd NAND3X1_327/A vdd NAND2X1
XNOR3X1_43 NOR3X1_43/A NOR3X1_43/B NOR3X1_43/C gnd NOR3X1_43/Y vdd NOR3X1
XNAND2X1_358 AND2X2_94/B AND2X2_94/A gnd OAI21X1_415/C vdd NAND2X1
XNOR3X1_32 NOR3X1_32/A NOR3X1_32/B NOR3X1_32/C gnd NOR3X1_33/C vdd NOR3X1
XNAND2X1_369 INVX1_306/A AND2X2_87/Y gnd NAND2X1_370/B vdd NAND2X1
XNOR3X1_21 NOR3X1_21/A NOR3X1_21/B NOR3X1_21/C gnd NOR3X1_21/Y vdd NOR3X1
XNAND2X1_347 INVX1_291/A OAI21X1_295/Y gnd AOI22X1_41/B vdd NAND2X1
XNOR3X1_10 NOR3X1_10/A NOR3X1_10/B NOR3X1_9/Y gnd NOR3X1_11/C vdd NOR3X1
XNAND3X1_9 INVX1_59/A NAND3X1_9/B INVX1_35/Y gnd INVX1_62/A vdd NAND3X1
XOAI21X1_116 NOR3X1_7/A NOR3X1_7/C NOR3X1_7/B gnd AOI21X1_49/A vdd OAI21X1
XOAI21X1_105 NOR3X1_13/A NOR3X1_13/B NAND3X1_72/A gnd NAND3X1_77/C vdd OAI21X1
XOAI21X1_149 AOI22X1_18/Y AOI21X1_66/Y AOI21X1_65/Y gnd AOI22X1_19/D vdd OAI21X1
XOAI21X1_138 INVX1_16/Y INVX1_148/Y NOR2X1_74/B gnd AOI21X1_60/B vdd OAI21X1
XOAI21X1_127 OAI22X1_5/A OAI22X1_5/B OAI21X1_127/C gnd XOR2X1_9/A vdd OAI21X1
XBUFX2_3 cos_alpha[0] gnd BUFX2_3/Y vdd BUFX2
XNAND2X1_177 cos_alpha[4] vertices[6] gnd OAI22X1_7/B vdd NAND2X1
XNAND2X1_155 cos_gamma[9] INVX1_9/A gnd INVX1_193/A vdd NAND2X1
XNAND2X1_111 INVX1_155/A OR2X2_15/Y gnd NAND3X1_80/A vdd NAND2X1
XNAND2X1_100 OAI21X1_85/Y NAND3X1_68/B gnd XNOR2X1_17/A vdd NAND2X1
XNAND2X1_122 dy[7] dx[7] gnd INVX1_131/A vdd NAND2X1
XNAND2X1_133 AND2X2_39/B AND2X2_39/A gnd AOI21X1_76/C vdd NAND2X1
XNAND2X1_166 NAND3X1_98/Y NAND3X1_95/Y gnd NAND2X1_536/B vdd NAND2X1
XNAND2X1_144 BUFX2_12/Y vertices[6] gnd INVX1_154/A vdd NAND2X1
XNAND2X1_199 cos_gamma[9] INVX1_27/Y gnd OAI21X1_311/A vdd NAND2X1
XNAND2X1_188 INVX1_171/Y NAND3X1_204/Y gnd AOI21X1_99/B vdd NAND2X1
XAOI21X1_3 AOI21X1_3/A INVX1_48/Y NOR2X1_36/Y gnd INVX1_49/A vdd AOI21X1
XXNOR2X1_77 XOR2X1_50/A XOR2X1_50/B gnd XNOR2X1_77/Y vdd XNOR2X1
XXNOR2X1_66 XNOR2X1_66/A XNOR2X1_66/B gnd XOR2X1_45/A vdd XNOR2X1
XXNOR2X1_44 XOR2X1_30/A XOR2X1_30/B gnd XNOR2X1_44/Y vdd XNOR2X1
XXNOR2X1_55 XNOR2X1_55/A XOR2X1_41/Y gnd XNOR2X1_56/B vdd XNOR2X1
XINVX1_90 INVX1_90/A gnd OR2X2_12/B vdd INVX1
XXNOR2X1_33 XNOR2X1_33/A INVX1_218/Y gnd XOR2X1_15/A vdd XNOR2X1
XXNOR2X1_22 NOR2X1_89/Y INVX1_157/Y gnd XOR2X1_10/A vdd XNOR2X1
XXNOR2X1_11 XNOR2X1_11/A INVX1_42/Y gnd OR2X2_7/A vdd XNOR2X1
XBUFX2_10 cos_alpha[2] gnd INVX1_15/A vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd vertices_out[14] vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd vertices_out[3] vdd BUFX2
XNOR2X1_1 INVX1_1/Y INVX1_2/Y gnd INVX1_9/A vdd NOR2X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_33 OAI21X1_81/Y INVX1_96/A NOR2X1_61/Y gnd NOR2X1_71/A vdd AOI21X1
XAOI21X1_55 INVX1_119/A INVX1_121/A NOR2X1_71/Y gnd NOR2X1_84/B vdd AOI21X1
XAOI21X1_44 NAND3X1_95/Y NAND3X1_98/Y INVX1_8/Y gnd INVX1_142/A vdd AOI21X1
XAOI21X1_22 NAND3X1_43/Y NAND3X1_44/Y INVX1_100/A gnd NOR3X1_4/B vdd AOI21X1
XAOI21X1_77 AOI21X1_77/A INVX1_162/A INVX1_140/A gnd NOR3X1_16/B vdd AOI21X1
XAOI21X1_11 OAI21X1_44/Y OAI21X1_45/Y INVX1_74/A gnd NOR3X1_1/C vdd AOI21X1
XOAI21X1_6 INVX1_1/Y INVX1_16/Y OR2X2_3/A gnd OAI21X1_7/C vdd OAI21X1
XAOI21X1_99 AND2X2_48/B AOI21X1_99/B INVX1_184/Y gnd NOR3X1_20/B vdd AOI21X1
XAOI21X1_66 AOI21X1_66/A AOI21X1_66/B AOI21X1_66/C gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_88 AOI21X1_88/A AOI21X1_88/B INVX1_178/A gnd AOI21X1_88/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XOAI21X1_491 OAI21X1_491/A XNOR2X1_63/A OAI21X1_491/C gnd INVX1_375/A vdd OAI21X1
XOAI21X1_480 NOR2X1_173/B OAI21X1_480/B OAI21X1_480/C gnd XOR2X1_52/B vdd OAI21X1
XXOR2X1_9 XOR2X1_9/A XOR2X1_9/B gnd XOR2X1_9/Y vdd XOR2X1
XNAND3X1_519 NAND3X1_519/A NAND3X1_519/B XOR2X1_44/Y gnd NAND3X1_522/A vdd NAND3X1
XNAND3X1_508 cos_gamma[2] NAND3X1_508/B NAND3X1_508/C gnd XOR2X1_43/A vdd NAND3X1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XINVX1_330 OR2X2_35/Y gnd INVX1_330/Y vdd INVX1
XINVX1_341 INVX1_341/A gnd INVX1_341/Y vdd INVX1
XINVX1_374 cos_alpha[15] gnd INVX1_374/Y vdd INVX1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XDFFPOSX1_11 BUFX2_28/A clk XOR2X1_16/Y gnd vdd DFFPOSX1
XFILL_27_0_0 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XNAND3X1_349 INVX1_280/A INVX1_279/Y OAI21X1_329/C gnd NAND3X1_350/C vdd NAND3X1
XNAND3X1_338 cos_gamma[9] INVX1_18/A NOR2X1_131/Y gnd AND2X2_82/B vdd NAND3X1
XNAND3X1_327 NAND3X1_327/A INVX1_295/A AOI22X1_35/D gnd NAND3X1_330/C vdd NAND3X1
XNAND3X1_316 AND2X2_80/A OAI21X1_301/C OAI21X1_299/Y gnd INVX1_270/A vdd NAND3X1
XNAND3X1_305 AOI22X1_41/A NAND3X1_305/B OAI21X1_294/Y gnd AND2X2_64/A vdd NAND3X1
XFILL_18_0_0 gnd vdd FILL
XNAND2X1_518 NOR2X1_191/A XNOR2X1_67/Y gnd AOI22X1_58/D vdd NAND2X1
XNAND2X1_507 vertices[7] cos_alpha[8] gnd XOR2X1_46/B vdd NAND2X1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XNAND2X1_529 OAI22X1_13/Y AND2X2_108/A gnd NOR3X1_45/C vdd NAND2X1
XAOI21X1_197 OAI21X1_325/C NOR2X1_141/Y NOR2X1_158/Y gnd INVX1_312/A vdd AOI21X1
XAOI21X1_164 OAI21X1_269/C XOR2X1_17/B NOR2X1_140/Y gnd INVX1_278/A vdd AOI21X1
XAOI21X1_175 OAI21X1_342/Y NAND3X1_357/A OAI21X1_337/Y gnd NOR3X1_31/A vdd AOI21X1
XAOI21X1_186 OAI21X1_356/Y AND2X2_89/B INVX1_273/A gnd OAI21X1_359/A vdd AOI21X1
XAOI21X1_142 OAI21X1_288/Y NAND3X1_294/Y OAI21X1_331/B gnd OAI21X1_291/A vdd AOI21X1
XAOI21X1_153 NAND3X1_312/C NAND3X1_312/B INVX1_249/A gnd NOR3X1_25/C vdd AOI21X1
XAOI21X1_120 AOI21X1_92/C AOI21X1_92/A INVX1_213/Y gnd OAI21X1_238/C vdd AOI21X1
XAOI21X1_131 NAND3X1_240/C NAND3X1_240/B OAI21X1_237/C gnd OAI21X1_267/B vdd AOI21X1
XNAND3X1_113 NOR3X1_19/A NOR3X1_12/Y AOI22X1_16/D gnd INVX1_136/A vdd NAND3X1
XNAND3X1_102 cos_gamma[1] NOR2X1_73/Y OAI21X1_173/A gnd AOI21X1_45/B vdd NAND3X1
XNAND3X1_146 NAND3X1_99/C NAND3X1_151/B NAND3X1_151/C gnd NAND3X1_154/C vdd NAND3X1
XNAND3X1_157 BUFX2_5/Y INVX1_142/Y NAND3X1_457/B gnd AOI21X1_73/B vdd NAND3X1
XNAND3X1_168 NOR2X1_69/Y AOI21X1_78/B AOI21X1_78/A gnd AOI21X1_80/B vdd NAND3X1
XNAND3X1_135 OAI21X1_176/A AOI22X1_20/D AOI22X1_20/C gnd AOI21X1_84/A vdd NAND3X1
XNAND3X1_124 BUFX2_17/Y vertices[7] NAND3X1_124/C gnd AOI21X1_63/B vdd NAND3X1
XNAND3X1_179 AOI21X1_91/A AOI21X1_91/B XNOR2X1_27/Y gnd NAND3X1_185/A vdd NAND3X1
XFILL_20_2 gnd vdd FILL
XOAI21X1_309 INVX1_224/A AOI22X1_38/Y OAI21X1_366/C gnd OAI21X1_309/Y vdd OAI21X1
XFILL_13_1 gnd vdd FILL
XNAND2X1_304 AOI22X1_39/C AOI22X1_39/D gnd XNOR2X1_37/B vdd NAND2X1
XNAND2X1_337 vertices[6] cos_alpha[6] gnd OR2X2_32/B vdd NAND2X1
XNAND2X1_315 INVX1_268/Y OAI21X1_319/Y gnd AND2X2_84/B vdd NAND2X1
XNAND2X1_326 NAND3X1_342/Y NAND3X1_343/Y gnd NAND3X1_380/A vdd NAND2X1
XNAND2X1_348 OAI21X1_406/A AOI22X1_41/Y gnd NAND2X1_351/B vdd NAND2X1
XNAND2X1_359 cos_gamma[12] INVX1_27/Y gnd OAI21X1_475/A vdd NAND2X1
XNOR3X1_44 NOR3X1_44/A NOR3X1_44/B NOR3X1_44/C gnd NOR3X1_44/Y vdd NOR3X1
XNOR3X1_33 NOR3X1_33/A NOR3X1_33/B NOR3X1_33/C gnd NOR3X1_35/C vdd NOR3X1
XNOR3X1_11 INVX1_92/Y NOR3X1_11/B NOR3X1_11/C gnd NOR3X1_11/Y vdd NOR3X1
XNOR3X1_22 NOR3X1_22/A NOR3X1_22/B NOR3X1_22/C gnd NOR3X1_22/Y vdd NOR3X1
XOAI21X1_117 NOR3X1_9/B NOR3X1_9/C NOR3X1_9/A gnd AOI21X1_54/A vdd OAI21X1
XOAI21X1_128 NOR3X1_7/A NOR3X1_7/B AOI21X1_47/B gnd INVX1_163/A vdd OAI21X1
XOAI21X1_106 NOR3X1_14/A NOR3X1_14/B OAI21X1_97/Y gnd NAND3X1_80/C vdd OAI21X1
XOAI21X1_139 AOI21X1_60/Y AOI21X1_61/Y INVX1_150/A gnd OAI21X1_139/Y vdd OAI21X1
XBUFX2_4 cos_alpha[0] gnd BUFX2_4/Y vdd BUFX2
XNAND2X1_156 cos_gamma[7] INVX1_43/A gnd XNOR2X1_30/B vdd NAND2X1
XNAND2X1_189 dy[9] dx[9] gnd INVX1_186/A vdd NAND2X1
XNAND2X1_134 XOR2X1_8/B XOR2X1_8/A gnd NAND2X1_135/A vdd NAND2X1
XNAND2X1_123 AND2X2_27/B AND2X2_27/A gnd NOR3X1_7/B vdd NAND2X1
XNAND2X1_112 vertices[2] cos_alpha[5] gnd INVX1_126/A vdd NAND2X1
XNAND2X1_101 NOR2X1_69/A NOR2X1_69/B gnd NAND2X1_102/A vdd NAND2X1
XNAND2X1_167 cos_gamma[2] NAND2X1_536/B gnd INVX1_184/A vdd NAND2X1
XNAND2X1_145 BUFX2_4/Y vertices[8] gnd NAND3X1_124/C vdd NAND2X1
XNAND2X1_178 BUFX2_13/Y vertices[7] gnd INVX1_178/A vdd NAND2X1
XAOI21X1_4 NAND3X1_6/C INVX1_75/A INVX1_47/Y gnd NOR3X1_2/A vdd AOI21X1
XXNOR2X1_12 NOR2X1_38/Y INVX1_55/Y gnd XOR2X1_5/A vdd XNOR2X1
XXNOR2X1_23 XNOR2X1_23/A XNOR2X1_23/B gnd XNOR2X1_23/Y vdd XNOR2X1
XBUFX2_33 BUFX2_33/A gnd vertices_out[15] vdd BUFX2
XXNOR2X1_45 XNOR2X1_45/A INVX1_324/Y gnd XOR2X1_31/A vdd XNOR2X1
XXNOR2X1_67 XOR2X1_45/A XOR2X1_45/B gnd XNOR2X1_67/Y vdd XNOR2X1
XXNOR2X1_56 XNOR2X1_56/A XNOR2X1_56/B gnd XNOR2X1_57/A vdd XNOR2X1
XXNOR2X1_78 XNOR2X1_78/A XNOR2X1_78/B gnd OR2X2_59/B vdd XNOR2X1
XXNOR2X1_34 XOR2X1_20/A XOR2X1_20/B gnd XNOR2X1_34/Y vdd XNOR2X1
XINVX1_80 dz[5] gnd INVX1_80/Y vdd INVX1
XBUFX2_22 BUFX2_22/A gnd vertices_out[4] vdd BUFX2
XBUFX2_11 cos_alpha[2] gnd BUFX2_11/Y vdd BUFX2
XINVX1_91 cos_gamma[6] gnd INVX1_91/Y vdd INVX1
XNOR2X1_2 dy[0] dx[0] gnd NOR2X1_4/A vdd NOR2X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_34 NAND3X1_96/A NAND3X1_60/B NOR2X1_60/Y gnd NOR2X1_73/B vdd AOI21X1
XAOI21X1_23 OAI21X1_74/Y NAND3X1_46/B OAI21X1_97/A gnd NOR3X1_3/B vdd AOI21X1
XAOI21X1_12 NAND3X1_19/B NAND3X1_19/A OAI21X1_46/Y gnd OAI21X1_75/B vdd AOI21X1
XAOI21X1_45 AOI21X1_45/A AOI21X1_45/B INVX1_123/Y gnd NOR3X1_5/C vdd AOI21X1
XAOI21X1_56 NAND3X1_97/C NAND3X1_97/B NAND3X1_96/A gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_67 AND2X2_32/Y NAND3X1_82/C NOR3X1_14/Y gnd AOI21X1_67/Y vdd AOI21X1
XAOI21X1_78 AOI21X1_78/A AOI21X1_78/B NOR2X1_69/Y gnd NOR3X1_18/B vdd AOI21X1
XOAI21X1_7 OAI21X1_7/A OAI21X1_7/B OAI21X1_7/C gnd OAI21X1_8/C vdd OAI21X1
XAOI21X1_89 XNOR2X1_21/Y AOI22X1_18/D INVX1_181/Y gnd AOI21X1_89/Y vdd AOI21X1
XFILL_5_2_1 gnd vdd FILL
XFILL_13_1_1 gnd vdd FILL
XOAI21X1_481 INVX1_360/Y NOR2X1_177/A INVX1_361/A gnd INVX1_370/A vdd OAI21X1
XOAI21X1_492 INVX1_2/Y INVX1_374/Y INVX1_375/A gnd OAI21X1_492/Y vdd OAI21X1
XOAI21X1_470 OAI21X1_471/A OAI21X1_471/B AND2X2_103/Y gnd OAI21X1_470/Y vdd OAI21X1
XNAND3X1_509 cos_gamma[1] INVX1_370/Y NAND3X1_509/C gnd NAND3X1_510/A vdd NAND3X1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XINVX1_386 INVX1_386/A gnd INVX1_386/Y vdd INVX1
XINVX1_353 XOR2X1_36/Y gnd INVX1_353/Y vdd INVX1
XINVX1_331 INVX1_331/A gnd INVX1_331/Y vdd INVX1
XINVX1_320 INVX1_320/A gnd NOR3X1_36/C vdd INVX1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XINVX1_342 INVX1_342/A gnd INVX1_342/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_12 BUFX2_29/A clk XNOR2X1_37/Y gnd vdd DFFPOSX1
XFILL_27_0_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XNAND3X1_328 NAND3X1_330/B NAND3X1_330/C OAI21X1_305/C gnd AOI22X1_37/C vdd NAND3X1
XNAND3X1_339 cos_gamma[11] INVX1_27/Y INVX1_265/A gnd AND2X2_82/A vdd NAND3X1
XNAND3X1_306 OAI21X1_294/C NAND3X1_306/B NAND3X1_306/C gnd INVX1_291/A vdd NAND3X1
XNAND3X1_317 INVX1_238/Y NAND3X1_317/B AND2X2_72/B gnd AOI22X1_34/A vdd NAND3X1
XFILL_18_0_1 gnd vdd FILL
XNAND2X1_519 XNOR2X1_73/A XNOR2X1_75/Y gnd AOI22X1_58/B vdd NAND2X1
XNAND2X1_508 cos_alpha[6] vertices[9] gnd XNOR2X1_68/B vdd NAND2X1
XINVX1_194 cos_gamma[10] gnd OAI22X1_8/A vdd INVX1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XAOI21X1_121 OAI21X1_238/Y INVX1_247/A INVX1_214/Y gnd OAI21X1_240/A vdd AOI21X1
XAOI21X1_132 OAI21X1_232/Y NAND3X1_235/A OAI21X1_236/C gnd OAI21X1_271/A vdd AOI21X1
XAOI21X1_110 NAND3X1_185/A NAND3X1_185/B OAI21X1_192/C gnd OAI21X1_222/A vdd AOI21X1
XAOI21X1_198 NAND3X1_403/C NAND3X1_403/B INVX1_311/A gnd OAI21X1_388/B vdd AOI21X1
XAOI21X1_165 NAND3X1_346/C NAND3X1_346/B INVX1_309/A gnd INVX1_279/A vdd AOI21X1
XAOI21X1_187 OAI21X1_355/Y NAND3X1_368/B INVX1_273/Y gnd OAI21X1_359/B vdd AOI21X1
XAOI21X1_176 NAND3X1_295/C OAI21X1_287/Y NOR3X1_24/Y gnd NOR3X1_32/A vdd AOI21X1
XAOI21X1_154 NAND3X1_315/C NAND3X1_315/B XOR2X1_21/Y gnd OAI21X1_301/A vdd AOI21X1
XAOI21X1_143 NAND3X1_237/C OAI21X1_235/Y INVX1_246/Y gnd OAI21X1_291/C vdd AOI21X1
XNAND3X1_103 INVX1_123/Y AOI21X1_45/B AOI21X1_45/A gnd AOI21X1_46/A vdd NAND3X1
XNAND3X1_114 INVX1_143/A NAND3X1_114/B NAND3X1_114/C gnd AND2X2_39/A vdd NAND3X1
XNAND3X1_158 INVX1_160/A AOI21X1_73/B AOI21X1_73/A gnd AOI21X1_74/A vdd NAND3X1
XNAND3X1_169 INVX1_137/A AOI21X1_80/B AOI21X1_80/A gnd NAND3X1_169/Y vdd NAND3X1
XNAND3X1_147 NAND3X1_99/Y OAI21X1_219/A NAND3X1_154/C gnd AOI21X1_82/B vdd NAND3X1
XNAND3X1_136 INVX1_182/A AOI21X1_94/A AOI22X1_19/D gnd AOI21X1_84/B vdd NAND3X1
XNAND3X1_125 INVX1_154/A AOI21X1_63/A AOI21X1_63/B gnd AOI21X1_86/B vdd NAND3X1
XFILL_20_3 gnd vdd FILL
XFILL_13_2 gnd vdd FILL
XNAND2X1_338 vertices[5] cos_alpha[6] gnd OAI21X1_333/A vdd NAND2X1
XNAND2X1_316 INVX1_268/A AND2X2_72/Y gnd NAND3X1_340/C vdd NAND2X1
XNAND2X1_327 XOR2X1_21/B XOR2X1_21/A gnd AND2X2_80/B vdd NAND2X1
XNAND2X1_349 INVX1_239/A AND2X2_78/A gnd OAI21X1_353/A vdd NAND2X1
XNAND2X1_305 NAND3X1_276/A NAND3X1_276/B gnd INVX1_257/A vdd NAND2X1
XNOR3X1_45 NOR3X1_45/A NOR3X1_45/B NOR3X1_45/C gnd NOR3X1_46/C vdd NOR3X1
XNOR3X1_34 NOR3X1_34/A NOR3X1_34/B NOR3X1_34/C gnd NOR3X1_34/Y vdd NOR3X1
XNOR3X1_23 NOR3X1_23/A NOR3X1_23/B NOR3X1_23/C gnd NOR3X1_23/Y vdd NOR3X1
XNOR3X1_12 NOR3X1_12/A NOR3X1_12/B NOR3X1_12/C gnd NOR3X1_12/Y vdd NOR3X1
XOAI21X1_118 NOR3X1_8/A NOR3X1_8/C NOR3X1_8/B gnd AOI21X1_52/A vdd OAI21X1
XOAI21X1_107 NOR3X1_14/A NOR3X1_14/B NOR3X1_14/C gnd NAND3X1_82/C vdd OAI21X1
XOAI21X1_129 OAI21X1_91/C OR2X2_18/B OR2X2_14/Y gnd INVX1_143/A vdd OAI21X1
XBUFX2_5 cos_gamma[0] gnd BUFX2_5/Y vdd BUFX2
XNAND2X1_124 cos_gamma[8] INVX1_9/A gnd XOR2X1_9/B vdd NAND2X1
XNAND2X1_135 NAND2X1_135/A AOI21X1_48/B gnd INVX1_161/A vdd NAND2X1
XNAND2X1_102 NAND2X1_102/A NOR3X1_17/A gnd NOR3X1_9/A vdd NAND2X1
XNAND2X1_113 NOR2X1_77/A NOR2X1_77/B gnd NAND3X1_75/C vdd NAND2X1
XNAND2X1_146 AOI22X1_19/B AOI22X1_19/A gnd OAI21X1_176/A vdd NAND2X1
XNAND2X1_168 OAI21X1_219/A NOR2X1_107/A gnd NAND2X1_185/B vdd NAND2X1
XNAND2X1_157 OAI21X1_168/Y INVX1_170/Y gnd XNOR2X1_24/A vdd NAND2X1
XNAND2X1_179 AND2X2_43/Y AND2X2_44/Y gnd AOI21X1_87/A vdd NAND2X1
XNOR2X1_190 XOR2X1_49/B XNOR2X1_74/Y gnd OAI22X1_10/B vdd NOR2X1
XAOI21X1_5 NAND3X1_3/C INVX1_31/A INVX1_17/A gnd AOI21X1_5/Y vdd AOI21X1
XXNOR2X1_46 XNOR2X1_46/A INVX1_301/A gnd XNOR2X1_46/Y vdd XNOR2X1
XXNOR2X1_57 XNOR2X1_57/A XNOR2X1_57/B gnd INVX1_366/A vdd XNOR2X1
XXNOR2X1_35 XOR2X1_18/A XOR2X1_18/B gnd XNOR2X1_35/Y vdd XNOR2X1
XXNOR2X1_13 NOR2X1_51/Y INVX1_80/Y gnd XOR2X1_6/A vdd XNOR2X1
XXNOR2X1_24 XNOR2X1_24/A OAI22X1_5/Y gnd XNOR2X1_25/A vdd XNOR2X1
XXNOR2X1_68 XNOR2X1_68/A XNOR2X1_68/B gnd XOR2X1_46/A vdd XNOR2X1
XXNOR2X1_79 XNOR2X1_79/A XNOR2X1_79/B gnd XNOR2X1_81/A vdd XNOR2X1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XBUFX2_23 BUFX2_23/A gnd vertices_out[5] vdd BUFX2
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XBUFX2_12 cos_alpha[2] gnd BUFX2_12/Y vdd BUFX2
XNOR2X1_3 INVX1_4/Y INVX1_5/Y gnd NOR2X1_4/B vdd NOR2X1
XFILL_22_1_2 gnd vdd FILL
XAOI21X1_13 NAND3X1_6/C INVX1_47/Y INVX1_75/Y gnd OAI21X1_50/C vdd AOI21X1
XAOI21X1_46 AOI21X1_46/A AND2X2_36/A XOR2X1_8/Y gnd NOR3X1_6/B vdd AOI21X1
XAOI21X1_35 NAND3X1_57/B NAND3X1_57/A NAND3X1_57/C gnd NOR2X1_73/A vdd AOI21X1
XAOI21X1_68 OR2X2_10/A NAND3X1_88/C INVX1_156/Y gnd AOI21X1_68/Y vdd AOI21X1
XAOI21X1_24 NAND3X1_50/A NAND3X1_50/B OAI21X1_75/Y gnd OAI21X1_95/B vdd AOI21X1
XAOI21X1_57 NAND3X1_85/A NAND3X1_85/B OAI21X1_95/Y gnd AOI21X1_57/Y vdd AOI21X1
XOAI21X1_8 INVX1_2/Y INVX1_15/Y OAI21X1_8/C gnd AND2X2_5/A vdd OAI21X1
XAOI21X1_79 AOI21X1_79/A INVX1_165/A INVX1_164/A gnd NOR3X1_17/B vdd AOI21X1
XFILL_5_2_2 gnd vdd FILL
XOAI22X1_10 OAI22X1_10/A OAI22X1_10/B OAI22X1_12/B OAI22X1_12/A gnd OAI22X1_10/Y vdd
+ OAI22X1
XFILL_13_1_2 gnd vdd FILL
XOAI21X1_482 INVX1_356/A OAI21X1_482/B OAI21X1_482/C gnd OAI21X1_482/Y vdd OAI21X1
XOAI21X1_471 OAI21X1_471/A OAI21X1_471/B OAI21X1_471/C gnd OAI21X1_471/Y vdd OAI21X1
XOAI21X1_493 OAI22X1_11/B OAI22X1_11/A INVX1_373/Y gnd OAI21X1_493/Y vdd OAI21X1
XOAI21X1_460 OAI21X1_461/A OAI21X1_461/B XOR2X1_39/Y gnd AOI22X1_55/D vdd OAI21X1
XINVX1_310 cos_alpha[13] gnd INVX1_310/Y vdd INVX1
XINVX1_376 INVX1_376/A gnd INVX1_376/Y vdd INVX1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XINVX1_321 NOR3X1_37/A gnd INVX1_321/Y vdd INVX1
XINVX1_332 XOR2X1_33/Y gnd INVX1_332/Y vdd INVX1
XINVX1_365 INVX1_365/A gnd INVX1_365/Y vdd INVX1
XINVX1_343 INVX1_343/A gnd INVX1_343/Y vdd INVX1
XOAI21X1_290 OAI21X1_331/A NOR3X1_24/Y OAI21X1_331/B gnd OAI21X1_290/Y vdd OAI21X1
XAND2X2_90 OR2X2_40/A OR2X2_40/B gnd AND2X2_90/Y vdd AND2X2
XFILL_1_2 gnd vdd FILL
XDFFPOSX1_13 BUFX2_30/A clk NOR2X1_153/Y gnd vdd DFFPOSX1
XFILL_27_0_2 gnd vdd FILL
XFILL_2_0_2 gnd vdd FILL
XNAND3X1_329 INVX1_225/Y AOI22X1_37/C AOI22X1_37/D gnd NAND3X1_334/B vdd NAND3X1
XNAND3X1_307 NAND3X1_307/A INVX1_291/A OAI21X1_295/Y gnd AND2X2_78/A vdd NAND3X1
XNAND3X1_318 INVX1_238/A NAND3X1_318/B NAND3X1_318/C gnd AOI22X1_34/B vdd NAND3X1
XFILL_18_0_2 gnd vdd FILL
XNAND2X1_509 OAI21X1_488/Y NAND3X1_513/Y gnd XOR2X1_49/B vdd NAND2X1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XINVX1_151 NOR2X1_75/B gnd INVX1_151/Y vdd INVX1
XFILL_20_2_0 gnd vdd FILL
XAOI21X1_166 OR2X2_29/Y INVX1_281/A AND2X2_73/Y gnd OAI21X1_330/C vdd AOI21X1
XAOI21X1_144 OAI21X1_285/Y NAND3X1_294/A OAI21X1_288/C gnd OAI21X1_331/A vdd AOI21X1
XAOI21X1_133 OAI21X1_229/C XOR2X1_14/B NOR2X1_122/Y gnd INVX1_243/A vdd AOI21X1
XAOI21X1_100 NAND3X1_205/C NAND3X1_205/B INVX1_184/A gnd NOR3X1_20/C vdd AOI21X1
XAOI21X1_155 AND2X2_54/Y AOI22X1_28/D INVX1_253/Y gnd OAI21X1_303/C vdd AOI21X1
XAOI21X1_111 INVX1_147/Y INVX1_205/Y NOR2X1_96/Y gnd INVX1_207/A vdd AOI21X1
XAOI21X1_122 OAI21X1_237/Y NAND3X1_239/B INVX1_214/A gnd OAI21X1_240/B vdd AOI21X1
XAOI21X1_199 NAND3X1_402/C NAND3X1_402/B INVX1_311/Y gnd OAI21X1_388/A vdd AOI21X1
XAOI21X1_177 OAI21X1_389/C OAI21X1_344/Y AND2X2_74/Y gnd NOR3X1_32/B vdd AOI21X1
XAOI21X1_188 AND2X2_92/B NAND3X1_380/C NAND3X1_380/A gnd OAI21X1_361/A vdd AOI21X1
XNAND3X1_104 NOR2X1_72/Y AOI22X1_15/C AND2X2_36/B gnd AND2X2_36/A vdd NAND3X1
XNAND3X1_148 INVX1_173/A AOI21X1_71/Y OAI21X1_153/Y gnd NAND3X1_200/A vdd NAND3X1
XNAND3X1_137 AOI21X1_84/A AOI21X1_84/B AOI21X1_67/Y gnd AOI21X1_70/A vdd NAND3X1
XNAND3X1_115 INVX1_143/Y NAND3X1_115/B NAND3X1_115/C gnd AND2X2_39/B vdd NAND3X1
XNAND3X1_126 INVX1_154/Y AOI22X1_24/D AOI22X1_17/D gnd AOI21X1_86/A vdd NAND3X1
XNAND3X1_159 INVX1_160/Y AOI22X1_21/C AOI22X1_21/D gnd AOI21X1_74/B vdd NAND3X1
XFILL_11_2_0 gnd vdd FILL
XNOR3X1_35 NOR3X1_35/A NOR3X1_35/B NOR3X1_35/C gnd NOR3X1_35/Y vdd NOR3X1
XNAND2X1_339 vertices[6] cos_alpha[7] gnd OAI21X1_442/A vdd NAND2X1
XNAND2X1_306 cos_gamma[12] INVX1_9/A gnd NOR2X1_163/A vdd NAND2X1
XNAND2X1_317 INVX1_268/Y AND2X2_72/Y gnd NAND3X1_341/C vdd NAND2X1
XNAND2X1_328 AND2X2_80/B AND2X2_80/A gnd NAND3X1_378/A vdd NAND2X1
XNOR3X1_24 NOR3X1_24/A NOR3X1_24/B NOR3X1_24/C gnd NOR3X1_24/Y vdd NOR3X1
XNOR3X1_13 NOR3X1_13/A NOR3X1_13/B NOR3X1_13/C gnd NOR3X1_13/Y vdd NOR3X1
XNOR3X1_46 INVX1_7/Y NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_46/Y vdd NOR3X1
XNAND3X1_90 INVX1_125/A NAND3X1_93/A NAND3X1_93/C gnd NAND3X1_96/B vdd NAND3X1
XNOR2X1_90 INVX1_91/Y INVX1_18/Y gnd NOR2X1_90/Y vdd NOR2X1
XNAND3X1_490 INVX1_363/A NAND3X1_492/B NAND3X1_492/A gnd NAND3X1_497/A vdd NAND3X1
XOAI21X1_119 AOI21X1_50/Y INVX1_135/Y INVX1_134/Y gnd AOI21X1_51/A vdd OAI21X1
XOAI21X1_108 AOI22X1_14/Y AOI21X1_42/Y NAND3X1_85/C gnd NAND3X1_88/C vdd OAI21X1
XBUFX2_6 cos_gamma[0] gnd INVX1_7/A vdd BUFX2
XNAND2X1_125 NOR2X1_84/A NOR2X1_84/B gnd AND2X2_34/B vdd NAND2X1
XNAND2X1_114 cos_alpha[3] vertices[4] gnd NOR2X1_76/B vdd NAND2X1
XNAND2X1_103 cos_gamma[4] AND2X2_13/Y gnd OAI21X1_92/B vdd NAND2X1
XNAND2X1_1 BUFX2_5/Y INVX1_9/A gnd INVX1_3/A vdd NAND2X1
XNAND2X1_147 AOI22X1_20/B AOI22X1_20/A gnd AOI21X1_94/A vdd NAND2X1
XNAND2X1_158 OR2X2_17/B OR2X2_17/A gnd AND2X2_47/B vdd NAND2X1
XNAND2X1_169 NAND3X1_132/B AOI22X1_19/A gnd OR2X2_21/A vdd NAND2X1
XNAND2X1_136 vertices[2] cos_alpha[6] gnd INVX1_147/A vdd NAND2X1
XFILL_25_1_0 gnd vdd FILL
XNOR2X1_191 NOR2X1_191/A XNOR2X1_67/Y gnd OAI22X1_11/C vdd NOR2X1
XNOR2X1_180 INVX1_364/Y XOR2X1_33/A gnd INVX1_367/A vdd NOR2X1
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 AOI21X1_6/A INVX1_62/A INVX1_24/A gnd NOR2X1_42/A vdd AOI21X1
XXNOR2X1_58 INVX1_383/A INVX1_366/Y gnd OR2X2_54/A vdd XNOR2X1
XXNOR2X1_36 XNOR2X1_36/A INVX1_250/Y gnd XOR2X1_21/A vdd XNOR2X1
XXNOR2X1_47 XNOR2X1_47/A INVX1_333/Y gnd OR2X2_47/B vdd XNOR2X1
XXNOR2X1_69 XOR2X1_48/A XOR2X1_48/B gnd XNOR2X1_73/A vdd XNOR2X1
XXNOR2X1_14 NOR2X1_52/Y INVX1_63/A gnd XNOR2X1_14/Y vdd XNOR2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XFILL_8_2_0 gnd vdd FILL
XXNOR2X1_25 XNOR2X1_25/A INVX1_193/A gnd XNOR2X1_26/B vdd XNOR2X1
XFILL_16_1_0 gnd vdd FILL
XINVX1_71 cos_alpha[5] gnd INVX1_71/Y vdd INVX1
XBUFX2_24 BUFX2_24/A gnd vertices_out[6] vdd BUFX2
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XDFFPOSX1_1 BUFX2_18/A clk NOR2X1_6/Y gnd vdd DFFPOSX1
XINVX1_82 XOR2X1_6/Y gnd INVX1_82/Y vdd INVX1
XBUFX2_13 cos_alpha[2] gnd BUFX2_13/Y vdd BUFX2
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd OR2X2_1/A vdd NOR2X1
XAOI21X1_58 NAND3X1_81/B NAND3X1_81/A OAI21X1_97/Y gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_47 AOI21X1_47/A AOI21X1_47/B AND2X2_27/Y gnd NOR3X1_8/A vdd AOI21X1
XAOI21X1_14 OAI21X1_49/Y OAI21X1_75/C NAND3X1_20/B gnd OAI21X1_51/A vdd AOI21X1
XAOI21X1_25 INVX1_77/Y OAI21X1_50/Y INVX1_104/Y gnd OAI21X1_78/C vdd AOI21X1
XAOI21X1_36 NAND3X1_59/C OAI21X1_79/Y NAND3X1_59/A gnd NAND3X1_97/A vdd AOI21X1
XAOI21X1_69 AOI21X1_95/B INVX1_183/A INVX1_155/Y gnd AOI21X1_69/Y vdd AOI21X1
XOAI21X1_9 INVX1_7/Y INVX1_18/Y INVX1_11/Y gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_11 OAI22X1_11/A OAI22X1_11/B OAI22X1_11/C OAI22X1_11/D gnd OAI22X1_11/Y vdd
+ OAI22X1
XOAI21X1_450 INVX1_10/Y INVX1_319/Y OAI21X1_450/C gnd OAI21X1_451/C vdd OAI21X1
XOAI21X1_494 OAI22X1_10/A OAI22X1_10/B INVX1_373/A gnd OAI21X1_494/Y vdd OAI21X1
XOAI21X1_472 OAI21X1_472/A XOR2X1_32/B OAI21X1_472/C gnd NOR2X1_178/B vdd OAI21X1
XOAI21X1_483 INVX1_353/Y OAI21X1_483/B OR2X2_53/Y gnd XOR2X1_44/A vdd OAI21X1
XOAI21X1_461 OAI21X1_461/A OAI21X1_461/B INVX1_362/Y gnd AOI22X1_54/D vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XINVX1_300 XOR2X1_25/Y gnd INVX1_300/Y vdd INVX1
XOAI21X1_280 NOR2X1_125/Y NOR2X1_126/Y INVX1_244/A gnd OAI21X1_280/Y vdd OAI21X1
XOAI21X1_291 OAI21X1_291/A OAI21X1_291/B OAI21X1_291/C gnd OAI21X1_291/Y vdd OAI21X1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XINVX1_355 INVX1_355/A gnd NOR3X1_44/A vdd INVX1
XINVX1_366 INVX1_366/A gnd INVX1_366/Y vdd INVX1
XINVX1_322 INVX1_322/A gnd INVX1_322/Y vdd INVX1
XINVX1_377 INVX1_377/A gnd NOR3X1_45/A vdd INVX1
XAND2X2_91 AND2X2_91/A AND2X2_91/B gnd AND2X2_91/Y vdd AND2X2
XINVX1_333 INVX1_333/A gnd INVX1_333/Y vdd INVX1
XAND2X2_80 AND2X2_80/A AND2X2_80/B gnd AND2X2_80/Y vdd AND2X2
XINVX1_344 INVX1_344/A gnd INVX1_344/Y vdd INVX1
XFILL_29_1 gnd vdd FILL
XDFFPOSX1_14 BUFX2_31/A clk XOR2X1_32/Y gnd vdd DFFPOSX1
XNAND3X1_308 INVX1_239/A AND2X2_64/Y AOI22X1_41/D gnd NAND3X1_308/Y vdd NAND3X1
XNAND3X1_319 AND2X2_80/A OAI21X1_299/Y AND2X2_65/Y gnd AOI22X1_34/C vdd NAND3X1
XINVX1_130 dz[7] gnd INVX1_130/Y vdd INVX1
XINVX1_141 NOR2X1_85/Y gnd OR2X2_16/B vdd INVX1
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_174 cos_alpha[9] gnd NOR2X1_95/B vdd INVX1
XINVX1_196 INVX1_196/A gnd OR2X2_23/A vdd INVX1
XINVX1_185 dz[9] gnd INVX1_185/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XAOI21X1_178 OAI21X1_345/Y NAND3X1_359/B OAI21X1_331/Y gnd NOR3X1_33/B vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_189 NAND3X1_379/B NAND3X1_379/C NAND3X1_379/A gnd OAI21X1_361/B vdd AOI21X1
XAOI21X1_167 OR2X2_32/Y OAI21X1_333/C INVX1_283/A gnd NOR3X1_26/B vdd AOI21X1
XAOI21X1_134 OAI21X1_231/Y INVX1_209/Y NOR3X1_21/B gnd NOR3X1_23/A vdd AOI21X1
XAOI21X1_145 INVX1_214/Y OAI21X1_238/Y INVX1_247/Y gnd OAI21X1_292/C vdd AOI21X1
XAOI21X1_101 NAND3X1_208/C AND2X2_48/A XOR2X1_11/Y gnd OAI21X1_200/A vdd AOI21X1
XAOI21X1_156 AND2X2_55/Y AOI22X1_29/D INVX1_254/Y gnd OAI21X1_304/C vdd AOI21X1
XAOI21X1_112 NAND3X1_180/A NAND3X1_180/B OAI21X1_189/C gnd OAI21X1_227/A vdd AOI21X1
XAOI21X1_123 NAND2X1_242/B OAI21X1_241/Y INVX1_8/Y gnd AOI22X1_31/B vdd AOI21X1
XNAND3X1_105 XOR2X1_8/Y AND2X2_36/A AOI21X1_46/A gnd AOI21X1_48/B vdd NAND3X1
XNAND3X1_138 INVX1_155/A AOI21X1_70/B AOI21X1_70/A gnd NAND3X1_144/A vdd NAND3X1
XNAND3X1_149 NAND3X1_96/C AOI21X1_83/B AOI21X1_83/A gnd NAND3X1_150/C vdd NAND3X1
XNAND3X1_127 AOI21X1_86/B AOI21X1_86/A AOI21X1_64/Y gnd AOI21X1_66/B vdd NAND3X1
XNAND3X1_116 AOI21X1_61/A INVX1_145/Y AOI21X1_61/B gnd NAND3X1_120/C vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XNAND2X1_307 INVX1_263/A INVX1_262/Y gnd INVX1_329/A vdd NAND2X1
XNAND2X1_318 INVX1_268/A OAI21X1_319/Y gnd NAND3X1_341/B vdd NAND2X1
XNOR3X1_47 NOR3X1_47/A NOR3X1_47/B NOR3X1_47/C gnd NOR3X1_49/C vdd NOR3X1
XNOR3X1_36 NOR3X1_36/A XOR2X1_30/Y NOR3X1_36/C gnd NOR3X1_37/C vdd NOR3X1
XNAND2X1_329 cos_gamma[1] AOI22X1_45/B gnd OAI21X1_356/C vdd NAND2X1
XNOR3X1_25 NOR3X1_25/A NOR3X1_25/B NOR3X1_25/C gnd NOR3X1_25/Y vdd NOR3X1
XNOR3X1_14 NOR3X1_14/A NOR3X1_14/B NOR3X1_14/C gnd NOR3X1_14/Y vdd NOR3X1
XNAND3X1_91 NAND3X1_97/A NAND3X1_96/B NAND3X1_96/C gnd NAND3X1_99/C vdd NAND3X1
XNAND3X1_80 NAND3X1_80/A NAND3X1_80/B NAND3X1_80/C gnd NAND3X1_85/A vdd NAND3X1
XNOR2X1_91 NOR2X1_91/A NOR2X1_7/B gnd NOR2X1_91/Y vdd NOR2X1
XNOR2X1_80 NOR2X1_80/A NOR2X1_80/B gnd NOR2X1_80/Y vdd NOR2X1
XNAND3X1_491 NAND3X1_498/A NAND3X1_497/A OAI21X1_466/Y gnd AOI22X1_60/A vdd NAND3X1
XNAND3X1_480 BUFX2_8/Y NAND3X1_480/B NAND3X1_509/C gnd NAND3X1_483/B vdd NAND3X1
XBUFX2_7 cos_gamma[0] gnd BUFX2_7/Y vdd BUFX2
XOAI21X1_109 AOI22X1_14/Y AOI21X1_42/Y OAI21X1_95/Y gnd NAND3X1_89/B vdd OAI21X1
XNAND2X1_104 OAI21X1_93/Y OR2X2_14/Y gnd NOR2X1_71/B vdd NAND2X1
XNAND2X1_148 AOI21X1_82/B AOI21X1_82/A gnd NAND3X1_457/B vdd NAND2X1
XNAND2X1_126 cos_gamma[3] AND2X2_13/Y gnd OR2X2_18/B vdd NAND2X1
XNAND2X1_159 AND2X2_47/B OR2X2_17/Y gnd NAND3X1_214/B vdd NAND2X1
XNAND2X1_115 BUFX2_13/Y vertices[5] gnd INVX1_127/A vdd NAND2X1
XNAND2X1_137 INVX1_149/Y INVX1_147/Y gnd AOI21X1_60/A vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XNAND2X1_2 dz[0] OR2X2_1/A gnd AND2X2_1/B vdd NAND2X1
XNOR2X1_181 XOR2X1_35/B XOR2X1_35/A gnd NOR2X1_181/Y vdd NOR2X1
XNOR2X1_192 XOR2X1_45/Y NOR2X1_192/B gnd OAI22X1_11/D vdd NOR2X1
XNOR2X1_170 AND2X2_89/Y XOR2X1_26/Y gnd NOR2X1_170/Y vdd NOR2X1
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_7 NAND3X1_9/B INVX1_59/A INVX1_35/Y gnd AOI21X1_7/Y vdd AOI21X1
XXNOR2X1_48 XNOR2X1_48/A INVX1_349/Y gnd INVX1_356/A vdd XNOR2X1
XXNOR2X1_59 XOR2X1_52/A XOR2X1_52/B gnd XNOR2X1_59/Y vdd XNOR2X1
XINVX1_50 vertices[4] gnd INVX1_50/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XXNOR2X1_15 XNOR2X1_15/A INVX1_95/Y gnd OR2X2_9/B vdd XNOR2X1
XFILL_8_2_1 gnd vdd FILL
XXNOR2X1_26 XNOR2X1_26/A XNOR2X1_26/B gnd OR2X2_17/A vdd XNOR2X1
XXNOR2X1_37 XNOR2X1_37/A XNOR2X1_37/B gnd XNOR2X1_37/Y vdd XNOR2X1
XFILL_16_1_1 gnd vdd FILL
XBUFX2_25 BUFX2_25/A gnd vertices_out[7] vdd BUFX2
XDFFPOSX1_2 BUFX2_19/A clk NOR2X1_13/Y gnd vdd DFFPOSX1
XBUFX2_14 cos_alpha[1] gnd INVX1_10/A vdd BUFX2
XNOR2X1_5 INVX1_3/Y NOR2X1_5/B gnd NOR2X1_6/A vdd NOR2X1
XAOI21X1_48 AOI21X1_48/A AOI21X1_48/B AOI21X1_48/C gnd NOR3X1_7/A vdd AOI21X1
XAOI21X1_26 OAI21X1_77/Y OAI21X1_95/C NOR2X1_59/Y gnd OAI21X1_79/A vdd AOI21X1
XAOI21X1_37 OAI21X1_72/Y NAND3X1_45/B OAI21X1_74/C gnd OAI21X1_97/B vdd AOI21X1
XAOI21X1_15 NAND3X1_8/A NAND3X1_8/B NAND3X1_8/C gnd NOR2X1_48/B vdd AOI21X1
XAOI21X1_59 OAI21X1_98/Y INVX1_126/Y NOR2X1_76/Y gnd INVX1_150/A vdd AOI21X1
XOAI22X1_12 OAI22X1_12/A OAI22X1_12/B OAI22X1_12/C OAI22X1_12/D gnd OAI22X1_12/Y vdd
+ OAI22X1
XOAI21X1_462 OAI21X1_464/B AOI22X1_54/Y INVX1_347/Y gnd OAI21X1_462/Y vdd OAI21X1
XOAI21X1_473 INVX1_331/Y INVX1_332/Y OAI21X1_473/C gnd NOR3X1_52/A vdd OAI21X1
XOAI21X1_484 OAI21X1_484/A XNOR2X1_68/A OR2X2_51/Y gnd XNOR2X1_62/B vdd OAI21X1
XOAI21X1_440 OAI21X1_440/A INVX1_316/Y AND2X2_91/A gnd OR2X2_50/B vdd OAI21X1
XOAI21X1_451 OR2X2_40/B XNOR2X1_70/A OAI21X1_451/C gnd OR2X2_56/A vdd OAI21X1
XOAI21X1_495 OAI21X1_495/A OAI21X1_495/B XNOR2X1_76/Y gnd OAI21X1_495/Y vdd OAI21X1
XNAND2X1_490 cos_gamma[15] INVX1_9/A gnd XNOR2X1_57/B vdd NAND2X1
XFILL_5_0_1 gnd vdd FILL
XINVX1_312 INVX1_312/A gnd INVX1_312/Y vdd INVX1
XOAI21X1_270 NOR2X1_102/A NOR2X1_140/A XOR2X1_17/Y gnd OAI21X1_270/Y vdd OAI21X1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XINVX1_323 INVX1_323/A gnd INVX1_323/Y vdd INVX1
XOAI21X1_281 INVX1_10/Y OAI22X1_9/D NOR2X1_149/A gnd OAI21X1_281/Y vdd OAI21X1
XINVX1_334 INVX1_334/A gnd INVX1_334/Y vdd INVX1
XOAI21X1_292 OAI21X1_293/A OAI21X1_293/B OAI21X1_292/C gnd OAI21X1_292/Y vdd OAI21X1
XINVX1_356 INVX1_356/A gnd INVX1_356/Y vdd INVX1
XINVX1_367 INVX1_367/A gnd OR2X2_54/B vdd INVX1
XAND2X2_92 AND2X2_92/A AND2X2_92/B gnd AND2X2_92/Y vdd AND2X2
XAND2X2_81 AND2X2_84/A AND2X2_81/B gnd AND2X2_81/Y vdd AND2X2
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XAND2X2_70 OR2X2_30/Y AND2X2_70/B gnd AND2X2_71/A vdd AND2X2
XINVX1_345 INVX1_345/A gnd INVX1_345/Y vdd INVX1
XDFFPOSX1_15 BUFX2_32/A clk NOR2X1_179/Y gnd vdd DFFPOSX1
XNAND3X1_309 BUFX2_5/Y NOR2X1_137/A AOI22X1_45/B gnd NAND3X1_312/C vdd NAND3X1
XINVX1_153 vertices[8] gnd OAI22X1_6/D vdd INVX1
XINVX1_186 INVX1_186/A gnd NOR2X1_99/B vdd INVX1
XINVX1_131 INVX1_131/A gnd NOR2X1_80/B vdd INVX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd NOR3X1_16/A vdd INVX1
XINVX1_120 NOR2X1_70/Y gnd OR2X2_14/B vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XFILL_20_2_2 gnd vdd FILL
XAOI21X1_146 OAI21X1_291/Y INVX1_289/A XNOR2X1_35/Y gnd OAI21X1_293/A vdd AOI21X1
XAOI21X1_179 XNOR2X1_35/Y OAI21X1_291/Y INVX1_289/Y gnd NOR3X1_35/A vdd AOI21X1
XAOI21X1_168 OAI21X1_278/C XOR2X1_20/B NOR2X1_146/Y gnd NOR3X1_26/A vdd AOI21X1
XAOI21X1_135 OAI21X1_340/C OAI21X1_281/Y INVX1_244/Y gnd NOR3X1_23/B vdd AOI21X1
XAOI21X1_113 NAND3X1_232/A OAI21X1_230/Y INVX1_211/Y gnd OAI21X1_276/B vdd AOI21X1
XAOI21X1_102 OAI21X1_200/Y NAND3X1_211/B NAND3X1_211/A gnd OAI21X1_202/B vdd AOI21X1
XAOI21X1_157 INVX1_223/A OAI21X1_249/Y INVX1_255/Y gnd OAI21X1_306/C vdd AOI21X1
XAOI21X1_124 NAND3X1_261/C NAND3X1_261/B XOR2X1_15/Y gnd OAI21X1_246/A vdd AOI21X1
XNAND3X1_106 AOI21X1_48/C AOI21X1_48/B AOI21X1_48/A gnd AOI21X1_47/B vdd NAND3X1
XNAND3X1_139 AOI21X1_84/C AOI21X1_84/A AOI21X1_84/B gnd INVX1_183/A vdd NAND3X1
XNAND3X1_128 AOI21X1_66/B AOI21X1_66/A AOI21X1_66/C gnd AOI21X1_85/B vdd NAND3X1
XNAND3X1_117 NOR2X1_86/Y AOI21X1_60/B AOI21X1_60/A gnd OAI21X1_177/C vdd NAND3X1
XFILL_11_2_2 gnd vdd FILL
XNAND2X1_308 INVX1_263/Y INVX1_262/A gnd AOI22X1_43/B vdd NAND2X1
XNAND2X1_319 AND2X2_84/A AND2X2_81/B gnd NAND3X1_382/B vdd NAND2X1
XNOR3X1_48 NOR3X1_48/A NOR3X1_48/B NOR3X1_48/C gnd NOR3X1_48/Y vdd NOR3X1
XNOR3X1_37 NOR3X1_37/A NOR3X1_37/B NOR3X1_37/C gnd NOR3X1_38/C vdd NOR3X1
XNOR3X1_26 NOR3X1_26/A NOR3X1_26/B NOR3X1_26/C gnd NOR3X1_26/Y vdd NOR3X1
XNOR3X1_15 NOR3X1_15/A NOR3X1_15/B NOR3X1_15/C gnd NOR3X1_15/Y vdd NOR3X1
XNAND3X1_81 NAND3X1_81/A NAND3X1_81/B OAI21X1_97/Y gnd NAND3X1_82/B vdd NAND3X1
XNAND3X1_92 INVX1_125/A NAND3X1_92/B NAND3X1_92/C gnd NAND3X1_97/B vdd NAND3X1
XNAND3X1_70 INVX1_126/Y OAI21X1_98/Y NAND3X1_75/C gnd NAND3X1_70/Y vdd NAND3X1
XNOR2X1_81 NOR2X1_81/A NOR2X1_81/B gnd NOR2X1_81/Y vdd NOR2X1
XNOR2X1_70 INVX1_65/Y INVX1_18/Y gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_92 NOR2X1_92/A NOR2X1_92/B gnd NOR2X1_92/Y vdd NOR2X1
XNAND3X1_470 NAND3X1_470/A NAND3X1_470/B OAI21X1_497/B gnd NAND3X1_473/B vdd NAND3X1
XNAND3X1_492 NAND3X1_492/A NAND3X1_492/B INVX1_363/Y gnd NAND3X1_498/C vdd NAND3X1
XNAND3X1_481 OAI21X1_458/C NAND3X1_481/B NAND3X1_481/C gnd NAND3X1_507/B vdd NAND3X1
XBUFX2_8 cos_gamma[0] gnd BUFX2_8/Y vdd BUFX2
XNAND2X1_3 INVX1_3/Y NOR2X1_5/B gnd INVX1_6/A vdd NAND2X1
XNAND2X1_105 NOR2X1_71/A NOR2X1_71/B gnd INVX1_121/A vdd NAND2X1
XNAND2X1_149 INVX1_142/Y OAI21X1_218/A gnd AOI22X1_21/D vdd NAND2X1
XNAND2X1_116 BUFX2_17/Y vertices[6] gnd NOR2X1_78/A vdd NAND2X1
XNAND2X1_127 cos_gamma[4] NAND2X1_70/Y gnd OR2X2_19/B vdd NAND2X1
XNAND2X1_138 cos_alpha[4] vertices[5] gnd INVX1_152/A vdd NAND2X1
XFILL_25_1_2 gnd vdd FILL
XNOR2X1_160 OR2X2_40/A OR2X2_40/B gnd NOR2X1_160/Y vdd NOR2X1
XFILL_0_1_2 gnd vdd FILL
XNOR2X1_182 INVX1_45/Y INVX1_350/Y gnd NOR2X1_183/A vdd NOR2X1
XNOR2X1_171 OR2X2_47/B OR2X2_47/A gnd NOR2X1_171/Y vdd NOR2X1
XNOR2X1_193 XOR2X1_48/Y XOR2X1_49/Y gnd OAI22X1_11/A vdd NOR2X1
XAOI21X1_8 AOI21X1_8/A INVX1_88/A NOR2X1_29/Y gnd NOR2X1_41/A vdd AOI21X1
XXNOR2X1_49 OR2X2_50/A OR2X2_50/B gnd XNOR2X1_49/Y vdd XNOR2X1
XINVX1_73 vertices[5] gnd INVX1_73/Y vdd INVX1
XXNOR2X1_38 XOR2X1_22/A XOR2X1_22/B gnd XNOR2X1_38/Y vdd XNOR2X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XXNOR2X1_16 NOR2X1_63/Y INVX1_106/Y gnd XOR2X1_7/A vdd XNOR2X1
XBUFX2_26 BUFX2_26/A gnd vertices_out[8] vdd BUFX2
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XFILL_8_2_2 gnd vdd FILL
XBUFX2_15 cos_alpha[1] gnd BUFX2_15/Y vdd BUFX2
XXNOR2X1_27 OAI22X1_7/D OAI22X1_7/C gnd XNOR2X1_27/Y vdd XNOR2X1
XFILL_16_1_2 gnd vdd FILL
XDFFPOSX1_3 BUFX2_20/A clk NOR2X1_22/Y gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A INVX1_6/Y gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 NAND2X1_70/Y BUFX2_9/Y INVX1_68/Y gnd OAI21X1_54/B vdd AOI21X1
XAOI21X1_49 AOI21X1_49/A AOI21X1_49/B AOI21X1_49/C gnd NOR3X1_9/B vdd AOI21X1
XAOI21X1_27 NAND3X1_24/Y NAND3X1_22/Y NAND3X1_54/Y gnd NAND3X1_58/C vdd AOI21X1
XAOI21X1_38 INVX1_101/Y INVX1_100/Y NOR2X1_58/Y gnd NOR3X1_13/C vdd AOI21X1
XOAI22X1_13 OAI22X1_13/A OAI22X1_13/B OAI22X1_13/C OAI22X1_13/D gnd OAI22X1_13/Y vdd
+ OAI22X1
XOAI21X1_496 INVX1_352/Y XNOR2X1_49/Y OAI21X1_496/C gnd XOR2X1_50/B vdd OAI21X1
XOAI21X1_452 NOR3X1_44/B NOR3X1_44/C NOR3X1_44/A gnd OAI21X1_452/Y vdd OAI21X1
XOAI21X1_463 AOI22X1_55/Y OAI21X1_479/A INVX1_347/A gnd OAI21X1_463/Y vdd OAI21X1
XOAI21X1_430 INVX1_322/Y OAI21X1_430/B OAI21X1_430/C gnd INVX1_357/A vdd OAI21X1
XOAI21X1_441 NOR3X1_38/A NOR3X1_38/B OAI21X1_441/C gnd INVX1_354/A vdd OAI21X1
XOAI21X1_485 XNOR2X1_52/B XOR2X1_37/Y OAI21X1_485/C gnd XNOR2X1_62/A vdd OAI21X1
XOAI21X1_474 INVX1_365/Y XOR2X1_33/A OR2X2_43/Y gnd XNOR2X1_56/A vdd OAI21X1
XNAND2X1_480 NAND3X1_481/C OAI21X1_458/Y gnd NAND2X1_481/B vdd NAND2X1
XNAND2X1_491 cos_gamma[12] INVX1_43/A gnd XNOR2X1_54/A vdd NAND2X1
XOAI21X1_90 INVX1_95/Y XNOR2X1_15/A OR2X2_13/Y gnd INVX1_119/A vdd OAI21X1
XFILL_5_0_2 gnd vdd FILL
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XINVX1_324 dz[13] gnd INVX1_324/Y vdd INVX1
XINVX1_313 INVX1_313/A gnd INVX1_313/Y vdd INVX1
XINVX1_357 INVX1_357/A gnd INVX1_357/Y vdd INVX1
XINVX1_302 OR2X2_41/B gnd OR2X2_35/B vdd INVX1
XINVX1_346 INVX1_346/A gnd INVX1_346/Y vdd INVX1
XOAI21X1_260 NOR2X1_116/A INVX1_231/Y INVX1_232/Y gnd OAI21X1_260/Y vdd OAI21X1
XINVX1_335 OR2X2_45/Y gnd OR2X2_46/B vdd INVX1
XOAI21X1_293 OAI21X1_293/A OAI21X1_293/B OAI21X1_293/C gnd OAI21X1_293/Y vdd OAI21X1
XOAI21X1_282 INVX1_10/Y OAI22X1_9/D AND2X2_63/Y gnd OAI21X1_282/Y vdd OAI21X1
XOAI21X1_271 OAI21X1_271/A OAI21X1_271/B INVX1_246/A gnd OAI21X1_289/C vdd OAI21X1
XAND2X2_93 AND2X2_93/A AND2X2_93/B gnd AND2X2_93/Y vdd AND2X2
XINVX1_379 INVX1_379/A gnd INVX1_379/Y vdd INVX1
XAND2X2_82 AND2X2_82/A AND2X2_82/B gnd XOR2X1_25/A vdd AND2X2
XAND2X2_71 AND2X2_71/A AND2X2_71/B gnd AND2X2_71/Y vdd AND2X2
XAND2X2_60 AND2X2_60/A AND2X2_60/B gnd INVX1_232/A vdd AND2X2
XDFFPOSX1_16 BUFX2_33/A clk NAND2X1_546/Y gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_132 XOR2X1_8/Y gnd NOR3X1_5/A vdd INVX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_165 INVX1_165/A gnd NOR3X1_16/C vdd INVX1
XINVX1_187 XOR2X1_11/Y gnd NOR3X1_20/A vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XAOI21X1_114 OAI21X1_279/C OAI21X1_231/Y INVX1_209/Y gnd OAI21X1_234/A vdd AOI21X1
XAOI21X1_103 OAI21X1_201/Y NAND3X1_214/A NAND3X1_214/B gnd OAI21X1_203/B vdd AOI21X1
XAOI21X1_169 OR2X2_33/Y OAI21X1_334/Y INVX1_284/Y gnd OAI21X1_386/B vdd AOI21X1
XAOI21X1_147 NAND3X1_297/C OAI21X1_289/Y XOR2X1_18/Y gnd OAI21X1_293/B vdd AOI21X1
XAOI21X1_136 OAI21X1_282/Y OAI21X1_283/Y INVX1_244/A gnd NOR3X1_23/C vdd AOI21X1
XAOI21X1_125 OAI21X1_246/Y NAND3X1_264/A NAND3X1_264/B gnd OAI21X1_248/B vdd AOI21X1
XAOI21X1_158 OAI21X1_305/Y NAND3X1_331/B INVX1_225/A gnd OAI21X1_307/B vdd AOI21X1
XNAND3X1_107 AOI21X1_47/B AOI21X1_47/A AND2X2_27/Y gnd AOI21X1_49/B vdd NAND3X1
XNAND3X1_129 AOI21X1_86/B AOI21X1_86/A AOI21X1_86/C gnd INVX1_181/A vdd NAND3X1
XNAND3X1_118 NAND3X1_120/C OAI21X1_177/C INVX1_150/Y gnd NAND3X1_132/B vdd NAND3X1
XNAND2X1_309 AOI22X1_43/B INVX1_329/A gnd INVX1_264/A vdd NAND2X1
XNOR3X1_49 XOR2X1_52/Y NOR3X1_49/B NOR3X1_49/C gnd NOR3X1_50/C vdd NOR3X1
XNOR3X1_38 NOR3X1_38/A NOR3X1_38/B NOR3X1_38/C gnd NOR3X1_39/C vdd NOR3X1
XNOR3X1_27 NOR3X1_27/A NOR3X1_27/B NOR3X1_27/C gnd NOR3X1_28/C vdd NOR3X1
XNOR3X1_16 NOR3X1_16/A NOR3X1_16/B NOR3X1_16/C gnd NOR3X1_17/C vdd NOR3X1
XFILL_20_0_0 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_60 NOR2X1_60/A INVX1_78/Y gnd NOR2X1_60/Y vdd NOR2X1
XNAND3X1_60 NAND3X1_96/A NAND3X1_60/B NOR2X1_60/Y gnd NAND3X1_95/A vdd NAND3X1
XNAND3X1_93 NAND3X1_93/A INVX1_125/Y NAND3X1_93/C gnd NAND3X1_97/C vdd NAND3X1
XNAND3X1_82 AND2X2_32/Y NAND3X1_82/B NAND3X1_82/C gnd NAND3X1_85/B vdd NAND3X1
XNOR2X1_71 NOR2X1_71/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XNAND3X1_71 INVX1_127/Y NAND3X1_71/B NAND3X1_71/C gnd NAND3X1_76/A vdd NAND3X1
XNOR2X1_82 NOR2X1_82/A NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XNAND3X1_471 INVX1_355/A NAND3X1_473/B NAND3X1_473/C gnd OAI21X1_482/C vdd NAND3X1
XNAND3X1_493 OAI21X1_467/Y NAND3X1_498/C AND2X2_102/Y gnd NAND3X1_494/B vdd NAND3X1
XNAND3X1_482 BUFX2_9/Y NAND3X1_507/B NAND3X1_528/B gnd NAND3X1_482/Y vdd NAND3X1
XNAND3X1_460 INVX1_346/Y NAND3X1_460/B OAI21X1_429/Y gnd NAND3X1_460/Y vdd NAND3X1
XNOR2X1_93 INVX1_65/Y OAI22X1_8/B gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 cos_gamma[0] gnd BUFX2_9/Y vdd BUFX2
XNAND2X1_106 XOR2X1_7/B XOR2X1_7/A gnd AND2X2_33/B vdd NAND2X1
XNAND2X1_128 OAI21X1_133/Y AND2X2_35/Y gnd NAND3X1_114/B vdd NAND2X1
XNAND2X1_4 BUFX2_2/Y vertices[1] gnd OAI21X1_7/A vdd NAND2X1
XNAND2X1_117 BUFX2_3/Y vertices[7] gnd NOR2X1_78/B vdd NAND2X1
XNAND2X1_139 NOR2X1_77/B INVX1_152/Y gnd NAND3X1_122/C vdd NAND2X1
XNOR2X1_150 dy[12] dx[12] gnd NOR2X1_151/A vdd NOR2X1
XNOR2X1_161 dy[13] dx[13] gnd NOR2X1_162/A vdd NOR2X1
XNOR2X1_183 NOR2X1_183/A XNOR2X1_63/Y gnd NOR2X1_184/A vdd NOR2X1
XNOR2X1_194 XNOR2X1_73/A XNOR2X1_75/Y gnd OAI22X1_11/B vdd NOR2X1
XNOR2X1_172 INVX1_36/Y NOR2X1_197/B gnd INVX1_342/A vdd NOR2X1
XAOI21X1_9 INVX1_39/Y INVX1_58/A NOR2X1_40/A gnd INVX1_64/A vdd AOI21X1
XXNOR2X1_39 XNOR2X1_39/A INVX1_292/Y gnd XOR2X1_24/A vdd XNOR2X1
XXNOR2X1_17 XNOR2X1_17/A XNOR2X1_17/B gnd XNOR2X1_17/Y vdd XNOR2X1
XXNOR2X1_28 OAI22X1_7/D INVX1_180/Y gnd XNOR2X1_28/Y vdd XNOR2X1
XINVX1_41 cos_gamma[2] gnd INVX1_41/Y vdd INVX1
XBUFX2_27 BUFX2_27/A gnd vertices_out[9] vdd BUFX2
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XBUFX2_16 cos_alpha[1] gnd BUFX2_16/Y vdd BUFX2
XDFFPOSX1_4 BUFX2_21/A clk XNOR2X1_10/Y gnd vdd DFFPOSX1
XNOR2X1_7 INVX1_8/Y NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XNAND3X1_290 NAND3X1_294/A OAI21X1_288/C OAI21X1_285/Y gnd OAI21X1_331/C vdd NAND3X1
XAOI21X1_17 NAND3X1_28/C AND2X2_26/A OAI21X1_39/Y gnd INVX1_83/A vdd AOI21X1
XAOI21X1_28 NAND3X1_63/C OAI21X1_80/Y XOR2X1_7/Y gnd INVX1_108/A vdd AOI21X1
XAOI21X1_39 NAND3X1_73/Y NAND3X1_74/Y INVX1_127/A gnd NOR3X1_13/A vdd AOI21X1
XOAI21X1_475 OAI21X1_475/A XOR2X1_40/A OR2X2_42/Y gnd XOR2X1_41/B vdd OAI21X1
XOAI21X1_497 OAI21X1_497/A OAI21X1_497/B AOI22X1_53/D gnd XOR2X1_50/A vdd OAI21X1
XOAI21X1_453 NOR3X1_44/B NOR3X1_44/C INVX1_355/A gnd OAI21X1_453/Y vdd OAI21X1
XOAI21X1_431 NOR3X1_40/A NOR3X1_40/B OAI21X1_431/C gnd INVX1_355/A vdd OAI21X1
XOAI21X1_486 OAI21X1_486/A XNOR2X1_64/A OR2X2_49/Y gnd XNOR2X1_66/A vdd OAI21X1
XOAI21X1_464 AOI22X1_54/Y OAI21X1_464/B INVX1_347/A gnd OAI21X1_464/Y vdd OAI21X1
XOAI21X1_420 OAI21X1_475/A XOR2X1_40/A OAI21X1_420/C gnd OR2X2_42/A vdd OAI21X1
XOAI21X1_442 OAI21X1_442/A OAI21X1_484/A OR2X2_39/Y gnd XOR2X1_36/B vdd OAI21X1
XNAND2X1_481 NAND3X1_478/Y NAND2X1_481/B gnd NAND3X1_509/C vdd NAND2X1
XNAND2X1_470 BUFX2_17/Y vertices[14] gnd XNOR2X1_70/A vdd NAND2X1
XFILL_8_0_0 gnd vdd FILL
XNAND2X1_492 cos_gamma[14] INVX1_27/Y gnd XOR2X1_40/B vdd NAND2X1
XOAI21X1_80 NOR2X1_61/Y AND2X2_25/Y INVX1_96/Y gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 INVX1_22/Y OAI22X1_8/B OAI21X1_91/C gnd OAI21X1_92/C vdd OAI21X1
XOAI21X1_250 AOI22X1_29/Y OAI21X1_250/B OAI21X1_250/C gnd AOI22X1_30/D vdd OAI21X1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XINVX1_314 INVX1_314/A gnd INVX1_314/Y vdd INVX1
XINVX1_347 INVX1_347/A gnd INVX1_347/Y vdd INVX1
XINVX1_369 INVX1_369/A gnd OR2X2_55/B vdd INVX1
XINVX1_358 INVX1_358/A gnd INVX1_358/Y vdd INVX1
XAND2X2_83 INVX1_301/Y AND2X2_83/B gnd OR2X2_41/B vdd AND2X2
XINVX1_303 INVX1_303/A gnd INVX1_303/Y vdd INVX1
XINVX1_336 INVX1_336/A gnd INVX1_336/Y vdd INVX1
XOAI21X1_272 INVX1_73/Y INVX1_148/Y OAI21X1_272/C gnd OAI21X1_273/C vdd OAI21X1
XAND2X2_50 XOR2X1_13/A XOR2X1_13/B gnd AND2X2_50/Y vdd AND2X2
XOAI21X1_283 INVX1_1/Y OAI22X1_9/B AND2X2_52/Y gnd OAI21X1_283/Y vdd OAI21X1
XAND2X2_72 AND2X2_72/A AND2X2_72/B gnd AND2X2_72/Y vdd AND2X2
XOAI21X1_294 OAI21X1_295/A OAI21X1_295/B OAI21X1_294/C gnd OAI21X1_294/Y vdd OAI21X1
XOAI21X1_261 INVX1_199/A AND2X2_48/Y AND2X2_61/A gnd OAI21X1_261/Y vdd OAI21X1
XAND2X2_61 AND2X2_61/A AND2X2_61/B gnd AND2X2_61/Y vdd AND2X2
XAND2X2_94 AND2X2_94/A AND2X2_94/B gnd AND2X2_94/Y vdd AND2X2
XFILL_23_2_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_177 vertices[6] gnd INVX1_177/Y vdd INVX1
XINVX1_144 cos_alpha[8] gnd NOR2X1_86/B vdd INVX1
XINVX1_133 NOR3X1_9/A gnd INVX1_133/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd NOR2X1_64/B vdd INVX1
XINVX1_122 NOR2X1_71/Y gnd INVX1_122/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_166 NOR3X1_19/Y gnd INVX1_166/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XFILL_27_1 gnd vdd FILL
XAOI21X1_137 OAI21X1_280/Y NAND3X1_291/B OAI21X1_286/C gnd OAI21X1_337/B vdd AOI21X1
XAOI21X1_148 OAI21X1_292/Y INVX1_274/A INVX1_240/Y gnd OAI21X1_295/A vdd AOI21X1
XAOI21X1_104 OAI21X1_203/Y AND2X2_57/B NOR2X1_84/Y gnd NOR3X1_22/A vdd AOI21X1
XAOI21X1_126 OAI21X1_247/Y NAND3X1_267/B NAND3X1_267/A gnd OAI21X1_250/B vdd AOI21X1
XAOI21X1_115 XNOR2X1_28/Y AOI21X1_90/A INVX1_212/Y gnd OAI21X1_235/C vdd AOI21X1
XAOI21X1_159 AOI22X1_39/Y OAI21X1_308/Y OAI21X1_309/Y gnd AOI22X1_44/D vdd AOI21X1
XNAND3X1_108 AOI21X1_49/B AOI21X1_49/A AOI21X1_49/C gnd AOI21X1_52/B vdd NAND3X1
XNAND3X1_119 NOR2X1_75/B NAND3X1_132/B OAI21X1_139/Y gnd AOI22X1_19/A vdd NAND3X1
XNOR3X1_17 NOR3X1_17/A NOR3X1_17/B NOR3X1_17/C gnd NOR3X1_18/C vdd NOR3X1
XNOR3X1_39 NOR3X1_39/A NOR3X1_39/B NOR3X1_39/C gnd NOR3X1_40/C vdd NOR3X1
XNOR3X1_28 NOR3X1_28/A NOR3X1_28/B NOR3X1_28/C gnd NOR3X1_29/C vdd NOR3X1
XFILL_20_0_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 NAND3X1_50/A NAND3X1_50/B OAI21X1_75/Y gnd OAI21X1_95/C vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_61 OR2X2_11/B OR2X2_11/A gnd NOR2X1_61/Y vdd NOR2X1
XNAND3X1_94 NAND3X1_96/A NAND3X1_97/B NAND3X1_97/C gnd NAND3X1_99/B vdd NAND3X1
XNOR2X1_50 dy[5] dx[5] gnd NOR2X1_51/A vdd NOR2X1
XNAND3X1_83 NAND3X1_85/B OAI21X1_95/Y NAND3X1_85/A gnd INVX1_156/A vdd NAND3X1
XNAND3X1_61 INVX1_7/A NAND3X1_61/B NAND3X1_95/A gnd OR2X2_11/A vdd NAND3X1
XNOR2X1_72 INVX1_41/Y OAI22X1_8/D gnd NOR2X1_72/Y vdd NOR2X1
XNAND3X1_72 NAND3X1_72/A NAND3X1_76/A NAND3X1_76/C gnd NAND3X1_78/A vdd NAND3X1
XNOR2X1_94 OR2X2_20/B OR2X2_20/A gnd NOR2X1_94/Y vdd NOR2X1
XNOR2X1_83 NOR2X1_83/A INVX1_18/Y gnd NOR2X1_83/Y vdd NOR2X1
XNAND3X1_494 AOI22X1_60/A NAND3X1_494/B XNOR2X1_46/Y gnd AOI22X1_60/B vdd NAND3X1
XNAND3X1_472 INVX1_356/A OAI21X1_452/Y OAI21X1_482/C gnd NAND3X1_472/Y vdd NAND3X1
XNAND3X1_450 INVX1_329/A NAND3X1_450/B OAI21X1_415/Y gnd NAND3X1_453/B vdd NAND3X1
XNAND3X1_483 INVX1_348/Y NAND3X1_483/B NAND3X1_483/C gnd NAND3X1_487/B vdd NAND3X1
XNAND3X1_461 cos_gamma[1] NAND3X1_508/B NAND3X1_508/C gnd NAND3X1_480/B vdd NAND3X1
XNAND2X1_107 AND2X2_33/B INVX1_109/A gnd AOI21X1_48/C vdd NAND2X1
XNAND2X1_129 AND2X2_35/B OR2X2_16/Y gnd OAI21X1_169/A vdd NAND2X1
XNAND2X1_5 vertices[1] BUFX2_15/Y gnd OR2X2_3/A vdd NAND2X1
XNAND2X1_118 AND2X2_24/Y AND2X2_31/Y gnd NAND3X1_71/C vdd NAND2X1
XNOR2X1_151 NOR2X1_151/A INVX1_293/Y gnd XNOR2X1_39/A vdd NOR2X1
XNOR2X1_162 NOR2X1_162/A INVX1_325/Y gnd XNOR2X1_45/A vdd NOR2X1
XNOR2X1_184 NOR2X1_184/A NOR2X1_184/B gnd XOR2X1_45/B vdd NOR2X1
XNOR2X1_195 OR2X2_58/B OR2X2_58/A gnd OAI22X1_13/C vdd NOR2X1
XNOR2X1_140 NOR2X1_140/A XOR2X1_23/A gnd NOR2X1_140/Y vdd NOR2X1
XNOR2X1_173 NOR2X1_173/A NOR2X1_173/B gnd NOR2X1_173/Y vdd NOR2X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XXNOR2X1_29 NOR2X1_99/Y INVX1_185/Y gnd XOR2X1_11/A vdd XNOR2X1
XXNOR2X1_18 NOR2X1_80/Y INVX1_130/Y gnd XOR2X1_8/A vdd XNOR2X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd NOR3X1_2/C vdd INVX1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XDFFPOSX1_5 BUFX2_22/A clk NOR2X1_41/Y gnd vdd DFFPOSX1
XBUFX2_28 BUFX2_28/A gnd vertices_out[10] vdd BUFX2
XBUFX2_17 cos_alpha[1] gnd BUFX2_17/Y vdd BUFX2
XNOR2X1_8 dy[1] dx[1] gnd NOR2X1_8/Y vdd NOR2X1
XNAND3X1_280 OAI21X1_258/Y OAI21X1_259/Y OAI21X1_316/C gnd INVX1_231/A vdd NAND3X1
XNAND3X1_291 NOR3X1_23/A NAND3X1_291/B OAI21X1_280/Y gnd NAND3X1_291/Y vdd NAND3X1
XAOI21X1_29 NAND3X1_66/C INVX1_135/A INVX1_134/A gnd NOR2X1_64/A vdd AOI21X1
XAOI21X1_18 NAND3X1_30/C OAI21X1_57/Y INVX1_64/Y gnd INVX1_86/A vdd AOI21X1
XOAI21X1_432 INVX1_312/A OAI21X1_432/B OAI21X1_432/C gnd INVX1_352/A vdd OAI21X1
XOAI21X1_410 OAI21X1_410/A NOR3X1_42/Y INVX1_327/A gnd AOI22X1_47/D vdd OAI21X1
XOAI21X1_421 OR2X2_36/B OR2X2_36/A OAI21X1_421/C gnd INVX1_339/A vdd OAI21X1
XOAI21X1_465 AOI22X1_55/Y OAI21X1_479/A INVX1_347/Y gnd OAI21X1_465/Y vdd OAI21X1
XOAI21X1_454 OAI21X1_456/A OAI21X1_456/B INVX1_358/A gnd OAI21X1_454/Y vdd OAI21X1
XOAI21X1_487 OR2X2_52/B OR2X2_52/A OR2X2_57/Y gnd OAI21X1_488/C vdd OAI21X1
XOAI21X1_443 INVX1_148/Y OAI22X1_6/D OAI21X1_443/C gnd OAI21X1_444/C vdd OAI21X1
XOAI21X1_498 INVX1_344/A INVX1_343/A INVX1_345/A gnd INVX1_378/A vdd OAI21X1
XOAI21X1_476 OAI21X1_476/A XNOR2X1_80/A OR2X2_44/Y gnd XNOR2X1_55/A vdd OAI21X1
XNAND2X1_460 OR2X2_50/B OR2X2_50/A gnd OAI21X1_496/C vdd NAND2X1
XNAND2X1_471 XOR2X1_36/Y XOR2X1_38/Y gnd NAND3X1_468/B vdd NAND2X1
XNAND2X1_493 OAI21X1_477/Y OR2X2_54/Y gnd INVX1_368/A vdd NAND2X1
XNAND2X1_482 NAND3X1_478/C OAI21X1_458/Y gnd NAND3X1_528/B vdd NAND2X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 INVX1_8/Y OAI22X1_8/D OR2X2_11/A gnd OAI21X1_81/Y vdd OAI21X1
XOAI21X1_70 INVX1_29/Y INVX1_28/Y AND2X2_22/Y gnd OAI21X1_70/Y vdd OAI21X1
XOAI21X1_92 OR2X2_13/A OAI21X1_92/B OAI21X1_92/C gnd OR2X2_14/A vdd OAI21X1
XOAI21X1_273 NOR2X1_142/A OR2X2_32/A OAI21X1_273/C gnd XOR2X1_19/A vdd OAI21X1
XOAI21X1_251 AOI22X1_30/Y OAI21X1_252/B AND2X2_57/Y gnd OAI21X1_251/Y vdd OAI21X1
XOAI21X1_240 OAI21X1_240/A OAI21X1_240/B INVX1_215/A gnd OAI21X1_240/Y vdd OAI21X1
XOAI21X1_262 OR2X2_19/A OR2X2_31/B OAI21X1_262/C gnd INVX1_238/A vdd OAI21X1
XINVX1_315 NOR3X1_40/A gnd INVX1_315/Y vdd INVX1
XINVX1_348 INVX1_348/A gnd INVX1_348/Y vdd INVX1
XAND2X2_95 AND2X2_95/A AND2X2_95/B gnd NOR3X1_43/A vdd AND2X2
XINVX1_326 XOR2X1_31/Y gnd NOR3X1_42/A vdd INVX1
XINVX1_359 INVX1_359/A gnd INVX1_359/Y vdd INVX1
XAND2X2_84 AND2X2_84/A AND2X2_84/B gnd OR2X2_41/A vdd AND2X2
XINVX1_304 INVX1_304/A gnd INVX1_304/Y vdd INVX1
XINVX1_337 INVX1_337/A gnd INVX1_337/Y vdd INVX1
XAND2X2_73 XOR2X1_19/Y INVX1_243/Y gnd AND2X2_73/Y vdd AND2X2
XAND2X2_62 XOR2X1_19/A XOR2X1_19/B gnd AND2X2_62/Y vdd AND2X2
XOAI21X1_284 NOR3X1_23/B NOR3X1_23/C NOR3X1_23/A gnd OAI21X1_284/Y vdd OAI21X1
XAND2X2_51 INVX1_208/A AND2X2_51/B gnd NOR3X1_21/C vdd AND2X2
XOAI21X1_295 OAI21X1_295/A OAI21X1_295/B OAI21X1_295/C gnd OAI21X1_295/Y vdd OAI21X1
XAND2X2_40 AND2X2_40/A AND2X2_40/B gnd OR2X2_20/B vdd AND2X2
XNAND2X1_290 cos_alpha[4] vertices[8] gnd AND2X2_75/A vdd NAND2X1
XFILL_23_2_2 gnd vdd FILL
XFILL_14_2_2 gnd vdd FILL
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_112 NOR3X1_12/A gnd INVX1_112/Y vdd INVX1
XINVX1_123 NOR2X1_72/Y gnd INVX1_123/Y vdd INVX1
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XINVX1_167 cos_gamma[8] gnd NOR2X1_91/A vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XINVX1_145 NOR2X1_86/Y gnd INVX1_145/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XFILL_27_2 gnd vdd FILL
XAOI21X1_149 OAI21X1_293/Y NAND3X1_302/B INVX1_240/A gnd OAI21X1_295/B vdd AOI21X1
XAOI21X1_138 OAI21X1_233/Y XNOR2X1_32/Y NOR2X1_106/Y gnd NOR3X1_24/C vdd AOI21X1
XAOI21X1_116 OAI21X1_276/C OAI21X1_233/Y XNOR2X1_32/Y gnd OAI21X1_236/B vdd AOI21X1
XAOI21X1_105 OAI21X1_205/Y NAND3X1_275/A NOR3X1_19/C gnd OAI21X1_308/B vdd AOI21X1
XAOI21X1_127 OAI21X1_249/Y INVX1_255/A INVX1_223/A gnd OAI21X1_252/B vdd AOI21X1
XNAND3X1_109 INVX1_133/Y AOI21X1_52/B AOI21X1_52/A gnd AOI21X1_54/B vdd NAND3X1
XNOR3X1_29 NOR3X1_29/A NOR3X1_29/B NOR3X1_29/C gnd NOR3X1_30/C vdd NOR3X1
XNOR3X1_18 NOR3X1_18/A NOR3X1_18/B NOR3X1_18/C gnd NOR3X1_19/C vdd NOR3X1
XFILL_20_0_2 gnd vdd FILL
XFILL_28_1_2 gnd vdd FILL
XFILL_3_1_2 gnd vdd FILL
XFILL_11_0_2 gnd vdd FILL
XNAND3X1_84 OR2X2_10/A INVX1_156/A NAND3X1_88/C gnd NAND3X1_92/B vdd NAND3X1
XNAND3X1_51 NOR2X1_59/Y OAI21X1_95/C OAI21X1_77/Y gnd INVX1_105/A vdd NAND3X1
XNAND3X1_40 INVX1_99/A OAI21X1_69/Y OAI21X1_70/Y gnd AOI22X1_9/B vdd NAND3X1
XNAND3X1_62 INVX1_96/A OAI21X1_81/Y OR2X2_11/Y gnd NAND3X1_63/C vdd NAND3X1
XNAND3X1_73 INVX1_1/A vertices[7] NOR2X1_78/A gnd NAND3X1_73/Y vdd NAND3X1
XFILL_19_1_2 gnd vdd FILL
XNOR2X1_73 NOR2X1_73/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XNOR2X1_51 NOR2X1_51/A INVX1_81/Y gnd NOR2X1_51/Y vdd NOR2X1
XNOR2X1_62 dy[6] dx[6] gnd NOR2X1_63/A vdd NOR2X1
XNOR2X1_40 NOR2X1_40/A INVX1_58/Y gnd NOR2X1_40/Y vdd NOR2X1
XNAND3X1_95 NAND3X1_95/A NAND3X1_99/B NAND3X1_99/C gnd NAND3X1_95/Y vdd NAND3X1
XNOR2X1_84 NOR2X1_84/A NOR2X1_84/B gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_95 INVX1_2/Y NOR2X1_95/B gnd OR2X2_21/B vdd NOR2X1
XNAND3X1_462 vertices[0] cos_alpha[14] INVX1_351/Y gnd OAI21X1_491/C vdd NAND3X1
XNAND3X1_473 NOR3X1_44/A NAND3X1_473/B NAND3X1_473/C gnd NAND3X1_476/C vdd NAND3X1
XNAND3X1_451 OAI21X1_415/C NAND3X1_451/B AND2X2_103/A gnd AND2X2_96/B vdd NAND3X1
XNAND3X1_495 INVX1_301/A NAND3X1_495/B NAND3X1_495/C gnd OAI21X1_473/C vdd NAND3X1
XNAND3X1_440 INVX1_340/A AOI22X1_46/D NAND3X1_440/C gnd NAND3X1_443/C vdd NAND3X1
XNAND3X1_484 BUFX2_5/Y NAND3X1_484/B NAND3X1_509/C gnd NAND3X1_485/B vdd NAND3X1
XNAND2X1_119 NAND3X1_70/Y OAI21X1_99/Y gnd NAND3X1_77/B vdd NAND2X1
XNAND2X1_108 vertices[1] cos_alpha[7] gnd NOR2X1_74/B vdd NAND2X1
XNAND2X1_6 dz[1] OR2X2_2/A gnd AND2X2_2/B vdd NAND2X1
XNOR2X1_185 XNOR2X1_67/Y NOR2X1_192/B gnd OAI22X1_12/A vdd NOR2X1
XNOR2X1_141 INVX1_45/Y INVX1_241/Y gnd NOR2X1_141/Y vdd NOR2X1
XNOR2X1_130 NOR2X1_163/A INVX1_260/Y gnd INVX1_261/A vdd NOR2X1
XNOR2X1_163 NOR2X1_163/A INVX1_299/Y gnd INVX1_365/A vdd NOR2X1
XNOR2X1_174 INVX1_41/Y NOR2X1_196/B gnd INVX1_348/A vdd NOR2X1
XNOR2X1_196 INVX1_22/Y NOR2X1_196/B gnd NOR2X1_196/Y vdd NOR2X1
XNOR2X1_152 NOR2X1_152/A NOR2X1_152/B gnd NOR2X1_153/B vdd NOR2X1
XXNOR2X1_19 NOR2X1_81/Y XNOR2X1_19/B gnd XNOR2X1_19/Y vdd XNOR2X1
XINVX1_32 dz[3] gnd INVX1_32/Y vdd INVX1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_54 NOR3X1_2/A gnd INVX1_54/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_65 cos_gamma[5] gnd INVX1_65/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XBUFX2_29 BUFX2_29/A gnd vertices_out[11] vdd BUFX2
XBUFX2_18 BUFX2_18/A gnd vertices_out[0] vdd BUFX2
XINVX1_98 INVX1_98/A gnd OR2X2_10/A vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XDFFPOSX1_6 BUFX2_23/A clk XNOR2X1_14/Y gnd vdd DFFPOSX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND3X1_292 OR2X2_29/Y INVX1_281/A OAI21X1_328/C gnd NAND3X1_292/Y vdd NAND3X1
XNAND3X1_281 INVX1_234/A AND2X2_67/B NAND3X1_324/C gnd AND2X2_67/A vdd NAND3X1
XAOI21X1_19 OAI21X1_55/Y INVX1_70/A INVX1_79/A gnd OR2X2_9/A vdd AOI21X1
XNAND3X1_270 OAI21X1_250/C NAND3X1_272/A NAND3X1_272/B gnd INVX1_255/A vdd NAND3X1
XOAI21X1_433 INVX1_16/Y INVX1_277/Y OR2X2_48/B gnd OAI21X1_434/C vdd OAI21X1
XOAI21X1_466 OAI21X1_467/A OAI21X1_467/B INVX1_363/Y gnd OAI21X1_466/Y vdd OAI21X1
XOAI21X1_455 OR2X2_58/A OAI21X1_457/B INVX1_358/Y gnd OAI21X1_455/Y vdd OAI21X1
XOAI21X1_411 AOI22X1_46/Y AOI22X1_47/Y OAI21X1_411/C gnd AOI22X1_49/D vdd OAI21X1
XOAI21X1_400 NOR3X1_37/B NOR3X1_37/C NOR3X1_37/A gnd OAI21X1_400/Y vdd OAI21X1
XOAI21X1_444 OAI21X1_484/A XNOR2X1_68/A OAI21X1_444/C gnd OR2X2_51/A vdd OAI21X1
XOAI21X1_422 OAI21X1_476/A XNOR2X1_80/A OAI22X1_8/Y gnd OR2X2_44/A vdd OAI21X1
XOAI21X1_477 INVX1_364/Y XOR2X1_33/A OR2X2_54/A gnd OAI21X1_477/Y vdd OAI21X1
XOAI21X1_488 NOR2X1_187/Y AND2X2_106/Y OAI21X1_488/C gnd OAI21X1_488/Y vdd OAI21X1
XOAI21X1_499 INVX1_36/Y OAI21X1_499/B NOR2X1_197/Y gnd OAI21X1_499/Y vdd OAI21X1
XNAND2X1_461 INVX1_352/Y XNOR2X1_49/Y gnd AOI22X1_53/B vdd NAND2X1
XNAND2X1_494 OR2X2_55/B OR2X2_55/A gnd AOI22X1_59/B vdd NAND2X1
XNAND2X1_472 OR2X2_53/B OR2X2_53/A gnd NAND2X1_473/A vdd NAND2X1
XNAND2X1_483 NAND3X1_484/B NAND3X1_482/Y gnd NAND3X1_483/C vdd NAND2X1
XNAND2X1_450 OAI21X1_428/C OAI21X1_478/A gnd NAND3X1_460/B vdd NAND2X1
XFILL_8_0_2 gnd vdd FILL
XFILL_8_1 gnd vdd FILL
XOAI21X1_82 INVX1_80/Y NOR2X1_51/A INVX1_81/A gnd XOR2X1_7/B vdd OAI21X1
XOAI21X1_60 INVX1_91/Y INVX1_9/Y NOR2X1_53/B gnd OAI21X1_60/Y vdd OAI21X1
XOAI21X1_93 INVX1_65/Y INVX1_18/Y OR2X2_14/A gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_71 INVX1_74/A AOI22X1_5/Y AOI22X1_3/D gnd OAI21X1_74/C vdd OAI21X1
XFILL_26_2_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XINVX1_316 INVX1_316/A gnd INVX1_316/Y vdd INVX1
XINVX1_305 INVX1_305/A gnd OR2X2_36/B vdd INVX1
XOAI21X1_274 OR2X2_34/A AND2X2_62/Y INVX1_243/A gnd INVX1_281/A vdd OAI21X1
XOAI21X1_285 OAI21X1_337/B NOR3X1_23/Y XOR2X1_20/Y gnd OAI21X1_285/Y vdd OAI21X1
XOAI21X1_296 INVX1_239/Y AOI22X1_32/Y OAI21X1_296/C gnd OAI21X1_296/Y vdd OAI21X1
XOAI21X1_230 NOR3X1_21/B NOR3X1_21/C NOR3X1_21/A gnd OAI21X1_230/Y vdd OAI21X1
XOAI21X1_263 OAI21X1_263/A OR2X2_37/B OAI21X1_263/C gnd OR2X2_28/A vdd OAI21X1
XOAI21X1_252 AOI22X1_30/Y OAI21X1_252/B AOI22X1_38/A gnd OAI21X1_252/Y vdd OAI21X1
XOAI21X1_241 OAI21X1_242/A NOR2X1_107/Y OAI21X1_354/B gnd OAI21X1_241/Y vdd OAI21X1
XINVX1_349 OR2X2_48/Y gnd INVX1_349/Y vdd INVX1
XAND2X2_96 AND2X2_96/A AND2X2_96/B gnd AND2X2_96/Y vdd AND2X2
XINVX1_327 INVX1_327/A gnd INVX1_327/Y vdd INVX1
XAND2X2_74 AND2X2_74/A AND2X2_74/B gnd AND2X2_74/Y vdd AND2X2
XINVX1_338 INVX1_338/A gnd INVX1_338/Y vdd INVX1
XAND2X2_85 AND2X2_97/B AND2X2_85/B gnd INVX1_304/A vdd AND2X2
XAND2X2_52 BUFX2_16/Y vertices[10] gnd AND2X2_52/Y vdd AND2X2
XAND2X2_63 BUFX2_3/Y vertices[11] gnd AND2X2_63/Y vdd AND2X2
XAND2X2_30 NOR2X1_78/A NOR2X1_78/B gnd AND2X2_30/Y vdd AND2X2
XAND2X2_41 OR2X2_20/A OR2X2_20/B gnd AND2X2_41/Y vdd AND2X2
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_291 BUFX2_11/Y vertices[9] gnd INVX1_244/A vdd NAND2X1
XNAND2X1_280 NAND3X1_202/C NAND2X1_280/B gnd AOI22X1_32/D vdd NAND2X1
XINVX1_146 cos_alpha[7] gnd INVX1_146/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_113 NOR3X1_12/B gnd INVX1_113/Y vdd INVX1
XINVX1_157 dz[8] gnd INVX1_157/Y vdd INVX1
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XINVX1_124 NOR2X1_73/Y gnd INVX1_124/Y vdd INVX1
XINVX1_168 NOR2X1_90/Y gnd INVX1_168/Y vdd INVX1
XINVX1_179 vertices[9] gnd OAI22X1_6/B vdd INVX1
XAOI21X1_139 OAI21X1_286/Y NAND3X1_291/Y XOR2X1_20/Y gnd NOR3X1_24/A vdd AOI21X1
XAOI21X1_117 OAI21X1_234/Y NAND3X1_232/Y XOR2X1_14/Y gnd OAI21X1_236/A vdd AOI21X1
XAOI21X1_106 NAND3X1_155/B NAND3X1_155/C NAND3X1_99/Y gnd NAND2X1_280/B vdd AOI21X1
XAOI21X1_128 XOR2X1_16/A XOR2X1_16/B INVX1_224/Y gnd XNOR2X1_37/A vdd AOI21X1
XFILL_23_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR3X1_19 NOR3X1_19/A NOR3X1_19/B NOR3X1_19/C gnd NOR3X1_19/Y vdd NOR3X1
XNAND3X1_96 NAND3X1_96/A NAND3X1_96/B NAND3X1_96/C gnd NAND3X1_98/B vdd NAND3X1
XNAND3X1_85 NAND3X1_85/A NAND3X1_85/B NAND3X1_85/C gnd NAND3X1_89/C vdd NAND3X1
XNAND3X1_52 INVX1_105/A OAI21X1_79/C OAI21X1_76/Y gnd INVX1_125/A vdd NAND3X1
XNAND3X1_63 XOR2X1_7/Y OAI21X1_80/Y NAND3X1_63/C gnd INVX1_109/A vdd NAND3X1
XNAND3X1_30 OAI21X1_57/Y INVX1_64/Y NAND3X1_30/C gnd INVX1_85/A vdd NAND3X1
XNAND3X1_41 INVX1_100/Y INVX1_101/Y AOI22X1_8/D gnd NAND3X1_45/B vdd NAND3X1
XNOR2X1_30 INVX1_36/Y NOR2X1_7/B gnd INVX1_37/A vdd NOR2X1
XNAND3X1_74 INVX1_10/A vertices[6] NOR2X1_78/B gnd NAND3X1_74/Y vdd NAND3X1
XNAND3X1_441 AND2X2_92/Y NAND3X1_443/B NAND3X1_443/C gnd AOI22X1_49/C vdd NAND3X1
XNAND3X1_430 INVX1_7/A NAND3X1_508/B NAND3X1_508/C gnd NOR2X1_173/B vdd NAND3X1
XNOR2X1_52 NOR2X1_52/A INVX1_89/Y gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_63 NOR2X1_63/A NOR2X1_63/B gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_41 NOR2X1_41/A INVX1_63/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_85 INVX1_65/Y INVX1_43/Y gnd NOR2X1_85/Y vdd NOR2X1
XNOR2X1_74 INVX1_97/A NOR2X1_74/B gnd NOR2X1_75/B vdd NOR2X1
XNOR2X1_96 OR2X2_22/B OR2X2_22/A gnd NOR2X1_96/Y vdd NOR2X1
XNAND3X1_463 INVX1_352/A OAI21X1_496/C OR2X2_50/Y gnd AOI22X1_53/A vdd NAND3X1
XNAND3X1_474 INVX1_356/Y OAI21X1_453/Y NAND3X1_476/C gnd NAND3X1_474/Y vdd NAND3X1
XNAND3X1_496 OAI21X1_471/C OAI21X1_469/Y AOI22X1_60/B gnd INVX1_385/A vdd NAND3X1
XNAND3X1_452 INVX1_329/Y AND2X2_96/B AOI22X1_52/D gnd AND2X2_96/A vdd NAND3X1
XNAND3X1_485 INVX1_348/A NAND3X1_485/B NAND3X1_485/C gnd OAI21X1_480/C vdd NAND3X1
XNAND2X1_7 OAI21X1_5/A XNOR2X1_1/Y gnd AND2X2_3/B vdd NAND2X1
XNAND2X1_109 vertices[3] cos_alpha[4] gnd NOR2X1_76/A vdd NAND2X1
XNOR2X1_142 NOR2X1_142/A OR2X2_32/A gnd OR2X2_34/B vdd NOR2X1
XNOR2X1_120 INVX1_205/A NOR2X1_142/A gnd OR2X2_29/B vdd NOR2X1
XNOR2X1_131 OAI22X1_8/A INVX1_43/Y gnd NOR2X1_131/Y vdd NOR2X1
XNOR2X1_186 NOR2X1_191/A XOR2X1_45/Y gnd OAI22X1_12/B vdd NOR2X1
XNOR2X1_175 NOR3X1_36/C NOR3X1_37/C gnd OR2X2_53/B vdd NOR2X1
XNOR2X1_164 XOR2X1_25/B XOR2X1_25/A gnd INVX1_364/A vdd NOR2X1
XNOR2X1_197 INVX1_65/Y NOR2X1_197/B gnd NOR2X1_197/Y vdd NOR2X1
XNOR2X1_153 NOR2X1_153/A NOR2X1_153/B gnd NOR2X1_153/Y vdd NOR2X1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_55 dz[4] gnd INVX1_55/Y vdd INVX1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_44 NOR3X1_2/B gnd INVX1_44/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_11 NOR2X1_7/Y gnd INVX1_11/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_22 cos_gamma[3] gnd INVX1_22/Y vdd INVX1
XDFFPOSX1_7 BUFX2_24/A clk XNOR2X1_17/Y gnd vdd DFFPOSX1
XBUFX2_19 BUFX2_19/A gnd vertices_out[1] vdd BUFX2
XNAND3X1_293 NOR2X1_121/Y OAI21X1_275/Y NAND3X1_293/C gnd NAND3X1_293/Y vdd NAND3X1
XNAND3X1_282 INVX1_234/Y NAND3X1_325/B NAND3X1_325/C gnd AOI22X1_35/B vdd NAND3X1
XNAND3X1_271 INVX1_223/A INVX1_255/A OAI21X1_249/Y gnd NAND3X1_276/A vdd NAND3X1
XNAND3X1_260 INVX1_217/Y AOI22X1_31/D NAND3X1_260/C gnd NAND3X1_261/C vdd NAND3X1
XOAI21X1_434 OAI21X1_491/A XNOR2X1_63/A OAI21X1_434/C gnd INVX1_351/A vdd OAI21X1
XOAI21X1_467 OAI21X1_467/A OAI21X1_467/B INVX1_363/A gnd OAI21X1_467/Y vdd OAI21X1
XOAI21X1_456 OAI21X1_456/A OAI21X1_456/B INVX1_358/Y gnd INVX1_377/A vdd OAI21X1
XOAI21X1_401 NOR3X1_39/B NOR3X1_39/C NOR3X1_39/A gnd OAI21X1_401/Y vdd OAI21X1
XOAI21X1_412 AOI22X1_46/Y AOI22X1_47/Y AND2X2_92/Y gnd AOI22X1_48/D vdd OAI21X1
XOAI21X1_478 OAI21X1_478/A AND2X2_100/Y OAI21X1_478/C gnd INVX1_369/A vdd OAI21X1
XOAI21X1_445 INVX1_177/Y NOR2X1_86/B OR2X2_51/A gnd OAI21X1_445/Y vdd OAI21X1
XOAI21X1_489 OR2X2_40/B XNOR2X1_70/A OR2X2_56/Y gnd XOR2X1_48/A vdd OAI21X1
XOAI21X1_423 INVX1_226/Y INVX1_43/Y OR2X2_44/A gnd AND2X2_98/B vdd OAI21X1
XNAND2X1_495 XOR2X1_39/B XOR2X1_39/A gnd NAND2X1_496/A vdd NAND2X1
XNAND2X1_473 NAND2X1_473/A OR2X2_53/Y gnd OAI21X1_483/B vdd NAND2X1
XNAND2X1_451 OAI21X1_478/C NAND3X1_460/Y gnd INVX1_347/A vdd NAND2X1
XNAND2X1_484 NAND3X1_480/B NAND3X1_482/Y gnd NAND3X1_485/C vdd NAND2X1
XNAND2X1_462 cos_alpha[7] vertices[8] gnd XNOR2X1_68/A vdd NAND2X1
XNAND2X1_440 cos_gamma[7] NAND3X1_457/B gnd XNOR2X1_79/A vdd NAND2X1
XOAI21X1_61 INVX1_69/A INVX1_83/A INVX1_84/A gnd INVX1_134/A vdd OAI21X1
XOAI21X1_50 OAI21X1_51/A INVX1_76/Y OAI21X1_50/C gnd OAI21X1_50/Y vdd OAI21X1
XOAI21X1_94 NOR2X1_71/Y INVX1_121/Y INVX1_119/Y gnd AND2X2_27/B vdd OAI21X1
XOAI21X1_83 INVX1_109/Y INVX1_108/A AND2X2_26/Y gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_72 INVX1_101/A NOR2X1_58/Y INVX1_100/A gnd OAI21X1_72/Y vdd OAI21X1
XFILL_26_2_1 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XINVX1_339 INVX1_339/A gnd INVX1_339/Y vdd INVX1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XINVX1_317 INVX1_317/A gnd INVX1_317/Y vdd INVX1
XOAI21X1_275 OR2X2_34/A AND2X2_62/Y INVX1_243/Y gnd OAI21X1_275/Y vdd OAI21X1
XOAI21X1_286 NOR3X1_23/B NOR3X1_23/C OAI21X1_286/C gnd OAI21X1_286/Y vdd OAI21X1
XOAI21X1_297 INVX1_239/Y AOI22X1_32/Y AND2X2_64/Y gnd OAI21X1_297/Y vdd OAI21X1
XOAI21X1_231 INVX1_1/Y OAI22X1_9/D INVX1_208/A gnd OAI21X1_231/Y vdd OAI21X1
XOAI21X1_264 INVX1_65/Y INVX1_124/Y OR2X2_28/A gnd OAI21X1_264/Y vdd OAI21X1
XOAI21X1_253 INVX1_193/A INVX1_195/Y OR2X2_27/A gnd AOI22X1_37/A vdd OAI21X1
XAND2X2_20 OR2X2_9/A OR2X2_9/B gnd AND2X2_20/Y vdd AND2X2
XOAI21X1_220 AOI21X1_97/C OAI21X1_220/B AOI21X1_96/B gnd INVX1_215/A vdd OAI21X1
XAND2X2_31 BUFX2_4/Y vertices[7] gnd AND2X2_31/Y vdd AND2X2
XOAI21X1_242 OAI21X1_242/A NOR2X1_107/Y OAI21X1_242/C gnd AOI22X1_41/D vdd OAI21X1
XAND2X2_97 AND2X2_97/A AND2X2_97/B gnd OR2X2_43/A vdd AND2X2
XAND2X2_86 AND2X2_86/A AND2X2_97/A gnd INVX1_305/A vdd AND2X2
XAND2X2_75 AND2X2_75/A AND2X2_75/B gnd AND2X2_75/Y vdd AND2X2
XNAND2X1_270 OAI21X1_264/Y OR2X2_28/Y gnd INVX1_236/A vdd NAND2X1
XAND2X2_64 AND2X2_64/A AND2X2_78/A gnd AND2X2_64/Y vdd AND2X2
XAND2X2_53 AND2X2_53/A AND2X2_53/B gnd AND2X2_53/Y vdd AND2X2
XAND2X2_42 OR2X2_22/A OR2X2_22/B gnd AND2X2_42/Y vdd AND2X2
XNAND2X1_281 vertices[2] cos_alpha[9] gnd OAI21X1_325/A vdd NAND2X1
XFILL_17_2_1 gnd vdd FILL
XNAND2X1_292 BUFX2_17/Y vertices[11] gnd NOR2X1_125/B vdd NAND2X1
XINVX1_114 cos_gamma[7] gnd NOR2X1_83/A vdd INVX1
XINVX1_169 NOR2X1_91/Y gnd NOR2X1_92/A vdd INVX1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd NOR2X1_89/B vdd INVX1
XINVX1_103 NOR2X1_58/A gnd INVX1_103/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd NOR2X1_81/B vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XAOI21X1_129 OAI21X1_316/C OAI21X1_259/Y OAI21X1_258/Y gnd NOR2X1_116/A vdd AOI21X1
XAOI21X1_118 OAI21X1_235/Y INVX1_246/A NAND3X1_237/C gnd OAI21X1_238/A vdd AOI21X1
XAOI21X1_107 INVX1_216/A NAND3X1_200/B AOI21X1_83/Y gnd OAI21X1_219/B vdd AOI21X1
XFILL_23_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XFILL_25_1 gnd vdd FILL
XNOR2X1_20 NOR2X1_20/A INVX1_20/Y gnd XNOR2X1_2/A vdd NOR2X1
XNAND3X1_97 NAND3X1_97/A NAND3X1_97/B NAND3X1_97/C gnd NAND3X1_98/C vdd NAND3X1
XNAND3X1_64 INVX1_109/A INVX1_108/Y OAI21X1_66/Y gnd INVX1_118/A vdd NAND3X1
XNAND3X1_86 INVX1_98/A NAND3X1_89/B NAND3X1_89/C gnd NAND3X1_92/C vdd NAND3X1
XNOR2X1_64 NOR2X1_64/A NOR2X1_64/B gnd NOR2X1_64/Y vdd NOR2X1
XNAND3X1_20 OAI21X1_75/C NAND3X1_20/B OAI21X1_49/Y gnd INVX1_76/A vdd NAND3X1
XNAND3X1_53 INVX1_125/A NAND3X1_59/A OAI21X1_78/Y gnd NAND3X1_57/A vdd NAND3X1
XNAND3X1_31 INVX1_38/A INVX1_85/A INVX1_86/Y gnd NAND3X1_32/B vdd NAND3X1
XNAND3X1_42 OAI21X1_74/C NAND3X1_45/B OAI21X1_72/Y gnd AOI22X1_9/C vdd NAND3X1
XNOR2X1_42 NOR2X1_42/A INVX1_60/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_31 XNOR2X1_5/B INVX1_67/A gnd NOR2X1_33/A vdd NOR2X1
XNAND3X1_75 INVX1_126/A OAI21X1_98/Y NAND3X1_75/C gnd NAND3X1_75/Y vdd NAND3X1
XNOR2X1_53 NOR2X1_82/A NOR2X1_53/B gnd INVX1_92/A vdd NOR2X1
XNAND3X1_475 INVX1_356/Y OAI21X1_452/Y OAI21X1_482/C gnd NAND3X1_475/Y vdd NAND3X1
XNAND3X1_453 NAND3X1_453/A NAND3X1_453/B AND2X2_96/A gnd OAI21X1_472/C vdd NAND3X1
XNAND3X1_442 NAND3X1_442/A AOI22X1_49/C AOI22X1_49/D gnd NAND3X1_446/A vdd NAND3X1
XNAND3X1_420 OAI21X1_379/Y NAND3X1_424/B OAI21X1_404/Y gnd INVX1_358/A vdd NAND3X1
XNAND3X1_464 cos_alpha[5] vertices[8] XOR2X1_30/A gnd OAI21X1_446/C vdd NAND3X1
XNAND3X1_431 INVX1_308/Y NAND3X1_431/B NAND3X1_431/C gnd NAND3X1_434/B vdd NAND3X1
XNOR2X1_75 NOR2X1_75/A NOR2X1_75/B gnd OR2X2_15/B vdd NOR2X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_86 INVX1_2/Y NOR2X1_86/B gnd NOR2X1_86/Y vdd NOR2X1
XNAND3X1_497 NAND3X1_497/A OAI21X1_466/Y AND2X2_102/Y gnd NAND3X1_497/Y vdd NAND3X1
XNAND3X1_486 INVX1_362/Y NAND3X1_487/B OAI21X1_480/C gnd AOI22X1_55/C vdd NAND3X1
XNAND2X1_8 XNOR2X1_1/B AND2X2_2/Y gnd OAI21X1_5/C vdd NAND2X1
XNOR2X1_176 dy[14] dx[14] gnd NOR2X1_177/A vdd NOR2X1
XNOR2X1_165 INVX1_365/A INVX1_364/A gnd XOR2X1_33/B vdd NOR2X1
XNOR2X1_143 OR2X2_34/B OR2X2_34/A gnd NOR2X1_143/Y vdd NOR2X1
XNOR2X1_154 INVX1_298/Y NOR2X1_7/B gnd INVX1_299/A vdd NOR2X1
XNOR2X1_121 OR2X2_29/B OR2X2_29/A gnd NOR2X1_121/Y vdd NOR2X1
XNOR2X1_110 NOR2X1_91/A INVX1_43/Y gnd INVX1_230/A vdd NOR2X1
XNOR2X1_132 NOR2X1_91/A OAI22X1_8/B gnd OR2X2_30/B vdd NOR2X1
XNOR2X1_187 XOR2X1_46/B XOR2X1_46/A gnd NOR2X1_187/Y vdd NOR2X1
XNOR2X1_198 NOR2X1_198/A NOR2X1_198/B gnd NOR2X1_198/Y vdd NOR2X1
XINVX1_45 vertices[1] gnd INVX1_45/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_12 dy[1] gnd NOR2X1_9/A vdd INVX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_34 OR2X2_6/Y gnd INVX1_34/Y vdd INVX1
XDFFPOSX1_8 BUFX2_25/A clk XNOR2X1_19/Y gnd vdd DFFPOSX1
XNAND3X1_294 NAND3X1_294/A OAI21X1_285/Y NOR3X1_24/C gnd NAND3X1_294/Y vdd NAND3X1
XNAND3X1_272 NAND3X1_272/A NAND3X1_272/B AND2X2_56/Y gnd AOI22X1_30/C vdd NAND3X1
XNAND3X1_250 INVX1_216/A AOI22X1_41/A NAND3X1_254/C gnd AOI22X1_32/A vdd NAND3X1
XNAND3X1_261 XOR2X1_15/Y NAND3X1_261/B NAND3X1_261/C gnd INVX1_222/A vdd NAND3X1
XNAND3X1_283 INVX1_238/A NAND3X1_317/B AND2X2_72/B gnd AND2X2_72/A vdd NAND3X1
XOAI21X1_435 INVX1_2/Y INVX1_350/Y INVX1_351/A gnd OAI21X1_435/Y vdd OAI21X1
XOAI21X1_479 OAI21X1_479/A INVX1_347/A OAI21X1_479/C gnd OR2X2_55/A vdd OAI21X1
XOAI21X1_402 NOR3X1_40/B NOR3X1_40/C NOR3X1_40/A gnd OAI21X1_402/Y vdd OAI21X1
XOAI21X1_457 OR2X2_58/A OAI21X1_457/B INVX1_358/A gnd OAI21X1_457/Y vdd OAI21X1
XOAI21X1_413 AOI22X1_48/Y AOI22X1_49/Y AND2X2_93/Y gnd AOI22X1_50/D vdd OAI21X1
XOAI21X1_468 INVX1_261/Y INVX1_300/Y XNOR2X1_46/A gnd OAI21X1_468/Y vdd OAI21X1
XOAI21X1_446 XOR2X1_29/A OR2X2_57/A OAI21X1_446/C gnd XNOR2X1_50/A vdd OAI21X1
XOAI21X1_424 INVX1_338/A INVX1_337/Y INVX1_336/Y gnd OAI21X1_424/Y vdd OAI21X1
XNAND2X1_452 XOR2X1_31/B XOR2X1_31/A gnd AOI22X1_55/A vdd NAND2X1
XNAND2X1_463 vertices[6] cos_alpha[8] gnd OR2X2_51/B vdd NAND2X1
XNAND2X1_430 NAND2X1_430/A OR2X2_43/Y gnd XOR2X1_33/A vdd NAND2X1
XNAND2X1_441 OAI21X1_424/Y NAND3X1_455/Y gnd OR2X2_46/A vdd NAND2X1
XNAND2X1_485 dy[14] dx[14] gnd INVX1_361/A vdd NAND2X1
XNAND2X1_496 NAND2X1_496/A AOI22X1_54/C gnd XOR2X1_52/A vdd NAND2X1
XNAND2X1_474 INVX1_353/Y OAI21X1_483/B gnd NAND3X1_468/C vdd NAND2X1
XOAI21X1_40 INVX1_47/A OAI21X1_40/B INVX1_75/A gnd OAI21X1_51/C vdd OAI21X1
XOAI21X1_73 NOR3X1_4/B NOR3X1_4/C NOR3X1_4/A gnd AOI22X1_9/D vdd OAI21X1
XOAI21X1_84 NOR2X1_64/A NOR2X1_64/B INVX1_93/A gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_95 OR2X2_10/Y OAI21X1_95/B OAI21X1_95/C gnd OAI21X1_95/Y vdd OAI21X1
XOAI21X1_51 OAI21X1_51/A INVX1_76/Y OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_62 INVX1_37/Y OAI21X1_64/A OAI21X1_62/C gnd INVX1_94/A vdd OAI21X1
XFILL_26_2_2 gnd vdd FILL
XFILL_1_2_2 gnd vdd FILL
XOAI21X1_221 INVX1_2/Y INVX1_203/Y NOR2X1_140/A gnd AND2X2_49/B vdd OAI21X1
XOAI21X1_210 INVX1_193/A INVX1_195/Y OAI21X1_210/C gnd OR2X2_24/B vdd OAI21X1
XINVX1_329 INVX1_329/A gnd INVX1_329/Y vdd INVX1
XINVX1_307 INVX1_307/A gnd INVX1_307/Y vdd INVX1
XINVX1_318 INVX1_318/A gnd INVX1_318/Y vdd INVX1
XOAI21X1_287 NOR3X1_24/A NOR3X1_24/B NOR3X1_24/C gnd OAI21X1_287/Y vdd OAI21X1
XOAI21X1_276 XOR2X1_14/Y OAI21X1_276/B OAI21X1_276/C gnd OAI21X1_288/C vdd OAI21X1
XOAI21X1_232 OAI21X1_276/B NOR2X1_106/Y XOR2X1_14/Y gnd OAI21X1_232/Y vdd OAI21X1
XOAI21X1_254 OR2X2_24/B OR2X2_24/A OR2X2_23/Y gnd INVX1_234/A vdd OAI21X1
XAND2X2_32 OR2X2_15/Y INVX1_155/A gnd AND2X2_32/Y vdd AND2X2
XOAI21X1_298 INVX1_218/Y NOR2X1_109/A INVX1_219/A gnd XOR2X1_21/B vdd OAI21X1
XAND2X2_21 AND2X2_21/A AND2X2_21/B gnd INVX1_110/A vdd AND2X2
XAND2X2_10 NAND3X1_8/C NAND3X1_3/Y gnd INVX1_43/A vdd AND2X2
XAND2X2_54 AND2X2_61/A AND2X2_54/B gnd AND2X2_54/Y vdd AND2X2
XOAI21X1_243 INVX1_7/Y NOR2X1_197/B OAI21X1_243/C gnd AOI22X1_31/D vdd OAI21X1
XOAI21X1_265 INVX1_220/Y OAI21X1_265/B AND2X2_65/B gnd OAI21X1_301/C vdd OAI21X1
XAND2X2_65 INVX1_222/A AND2X2_65/B gnd AND2X2_65/Y vdd AND2X2
XAND2X2_43 INVX1_10/A vertices[8] gnd AND2X2_43/Y vdd AND2X2
XNAND2X1_282 vertices[2] cos_alpha[10] gnd XOR2X1_23/A vdd NAND2X1
XNAND2X1_260 OAI21X1_260/Y NAND2X1_260/B gnd INVX1_233/A vdd NAND2X1
XAND2X2_98 OR2X2_44/Y AND2X2_98/B gnd INVX1_333/A vdd AND2X2
XAND2X2_87 AND2X2_87/A AND2X2_87/B gnd AND2X2_87/Y vdd AND2X2
XNAND2X1_293 AND2X2_52/Y AND2X2_63/Y gnd OAI21X1_340/C vdd NAND2X1
XAND2X2_76 BUFX2_15/Y vertices[12] gnd AND2X2_76/Y vdd AND2X2
XNAND2X1_271 INVX1_236/Y INVX1_237/Y gnd AND2X2_72/B vdd NAND2X1
XFILL_17_2_2 gnd vdd FILL
XINVX1_148 cos_alpha[6] gnd INVX1_148/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XINVX1_159 XOR2X1_10/Y gnd NOR3X1_15/A vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd NOR3X1_18/A vdd INVX1
XINVX1_115 NOR2X1_67/Y gnd NOR2X1_82/B vdd INVX1
XAOI21X1_119 OAI21X1_236/Y NAND3X1_236/A OAI21X1_271/B gnd OAI21X1_238/B vdd AOI21X1
XAOI21X1_108 NAND2X1_280/B NAND3X1_202/C OAI21X1_242/A gnd OAI21X1_354/A vdd AOI21X1
XFILL_23_0_2 gnd vdd FILL
XFILL_6_1_2 gnd vdd FILL
XFILL_14_0_2 gnd vdd FILL
XFILL_18_1 gnd vdd FILL
XNAND3X1_21 INVX1_76/A OAI21X1_47/Y OAI21X1_51/C gnd INVX1_104/A vdd NAND3X1
XNAND3X1_32 INVX1_87/A NAND3X1_32/B OAI21X1_58/Y gnd NOR3X1_12/A vdd NAND3X1
XNAND3X1_10 INVX1_24/A INVX1_62/A AOI21X1_6/A gnd INVX1_60/A vdd NAND3X1
XNAND3X1_65 INVX1_110/A INVX1_118/A OAI21X1_83/Y gnd INVX1_135/A vdd NAND3X1
XNAND3X1_87 NAND3X1_92/B INVX1_125/Y NAND3X1_92/C gnd NAND3X1_96/C vdd NAND3X1
XNOR2X1_65 OR2X2_12/B OR2X2_12/A gnd NOR3X1_12/C vdd NOR2X1
XNOR2X1_10 NOR2X1_8/Y NOR2X1_9/Y gnd OR2X2_2/A vdd NOR2X1
XNAND3X1_54 INVX1_53/A INVX1_54/Y INVX1_44/Y gnd NAND3X1_54/Y vdd NAND3X1
XNAND3X1_98 NOR2X1_73/A NAND3X1_98/B NAND3X1_98/C gnd NAND3X1_98/Y vdd NAND3X1
XNOR2X1_21 AND2X2_4/Y XOR2X1_3/Y gnd NOR2X1_22/A vdd NOR2X1
XNOR2X1_32 XNOR2X1_6/B XNOR2X1_6/A gnd NOR2X1_33/B vdd NOR2X1
XNAND3X1_76 NAND3X1_76/A NOR3X1_13/C NAND3X1_76/C gnd NAND3X1_77/A vdd NAND3X1
XNOR2X1_43 NOR2X1_43/A INVX1_37/Y gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_76 NOR2X1_76/A NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_54 INVX1_65/Y NOR2X1_7/B gnd INVX1_95/A vdd NOR2X1
XNAND3X1_43 BUFX2_2/Y vertices[6] NOR2X1_58/A gnd NAND3X1_43/Y vdd NAND3X1
XNOR2X1_87 INVX1_29/Y INVX1_71/Y gnd NOR2X1_87/Y vdd NOR2X1
XNAND3X1_476 INVX1_356/A OAI21X1_453/Y NAND3X1_476/C gnd NAND3X1_476/Y vdd NAND3X1
XNAND3X1_465 INVX1_354/A NAND3X1_468/B NAND3X1_468/C gnd AOI22X1_53/D vdd NAND3X1
XNAND3X1_498 NAND3X1_498/A OAI21X1_467/Y NAND3X1_498/C gnd NAND3X1_498/Y vdd NAND3X1
XNAND3X1_454 OAI21X1_472/C OAI21X1_417/Y NOR2X1_153/A gnd AOI22X1_56/C vdd NAND3X1
XNAND3X1_487 XOR2X1_39/Y NAND3X1_487/B OAI21X1_480/C gnd AOI22X1_54/C vdd NAND3X1
XNAND3X1_421 INVX1_322/Y OAI21X1_430/C OAI21X1_403/Y gnd NAND3X1_425/B vdd NAND3X1
XNAND3X1_443 OAI21X1_411/C NAND3X1_443/B NAND3X1_443/C gnd AOI22X1_48/C vdd NAND3X1
XNAND3X1_432 BUFX2_7/Y NAND3X1_432/B NAND3X1_432/C gnd AOI22X1_45/C vdd NAND3X1
XNAND3X1_410 INVX1_318/A OAI21X1_397/Y OR2X2_40/Y gnd NAND3X1_411/B vdd NAND3X1
XNOR2X1_98 dy[9] dx[9] gnd NOR2X1_99/A vdd NOR2X1
XNAND2X1_9 cos_gamma[2] INVX1_9/A gnd XOR2X1_1/B vdd NAND2X1
XNOR2X1_177 NOR2X1_177/A INVX1_361/Y gnd XNOR2X1_53/A vdd NOR2X1
XNOR2X1_155 INVX1_261/Y INVX1_300/Y gnd INVX1_301/A vdd NOR2X1
XNOR2X1_144 INVX1_50/Y NOR2X1_86/B gnd INVX1_283/A vdd NOR2X1
XNOR2X1_188 INVX1_71/Y OAI22X1_9/D gnd XOR2X1_48/B vdd NOR2X1
XNOR2X1_199 INVX1_226/Y OAI22X1_8/B gnd XNOR2X1_80/B vdd NOR2X1
XNOR2X1_166 NOR2X1_166/A NOR2X1_166/B gnd OR2X2_45/B vdd NOR2X1
XNOR2X1_122 OAI22X1_7/B NOR2X1_146/A gnd NOR2X1_122/Y vdd NOR2X1
XNOR2X1_111 NOR2X1_83/A OAI22X1_8/B gnd NOR2X1_113/A vdd NOR2X1
XNOR2X1_133 NOR2X1_133/A NOR2X1_166/A gnd NOR2X1_134/A vdd NOR2X1
XNOR2X1_100 OAI22X1_8/A NOR2X1_7/B gnd INVX1_195/A vdd NOR2X1
XINVX1_13 dx[1] gnd NOR2X1_9/B vdd INVX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XINVX1_46 cos_alpha[4] gnd INVX1_46/Y vdd INVX1
XINVX1_57 XOR2X1_5/Y gnd OR2X2_7/B vdd INVX1
XDFFPOSX1_9 BUFX2_26/A clk XNOR2X1_23/Y gnd vdd DFFPOSX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XNAND3X1_295 OAI21X1_331/C OAI21X1_287/Y NAND3X1_295/C gnd NAND3X1_298/A vdd NAND3X1
XNAND3X1_273 INVX1_223/Y AOI22X1_30/C AOI22X1_30/D gnd NAND3X1_276/B vdd NAND3X1
XNAND3X1_251 INVX1_201/A NAND3X1_251/B NAND3X1_251/C gnd NAND3X1_255/B vdd NAND3X1
XNAND3X1_262 INVX1_221/A INVX1_222/A NAND3X1_263/C gnd INVX1_253/A vdd NAND3X1
XNAND3X1_240 OAI21X1_237/C NAND3X1_240/B NAND3X1_240/C gnd INVX1_247/A vdd NAND3X1
XNAND3X1_284 INVX1_238/Y NAND3X1_318/B NAND3X1_318/C gnd AOI22X1_33/B vdd NAND3X1
XOAI21X1_403 NOR3X1_41/B NOR3X1_41/C NOR3X1_41/A gnd OAI21X1_403/Y vdd OAI21X1
XOAI21X1_414 AOI22X1_48/Y AOI22X1_49/Y OAI21X1_414/C gnd AOI22X1_51/D vdd OAI21X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_469 OAI21X1_511/A OAI21X1_469/B OAI21X1_511/B gnd OAI21X1_469/Y vdd OAI21X1
XOAI21X1_436 XOR2X1_23/B OAI21X1_437/C OR2X2_38/Y gnd XOR2X1_34/A vdd OAI21X1
XOAI21X1_425 NOR2X1_171/Y AND2X2_99/Y INVX1_339/A gnd OAI21X1_425/Y vdd OAI21X1
XOAI21X1_458 OAI21X1_458/A OAI21X1_458/B OAI21X1_458/C gnd OAI21X1_458/Y vdd OAI21X1
XOAI21X1_447 OR2X2_57/A OR2X2_57/B OAI22X1_9/Y gnd OR2X2_52/A vdd OAI21X1
XNAND2X1_497 INVX1_370/A OAI21X1_480/B gnd NAND3X1_510/B vdd NAND2X1
XNAND2X1_475 INVX1_353/Y XOR2X1_38/Y gnd NAND3X1_469/B vdd NAND2X1
XNAND2X1_486 OAI21X1_473/C OAI21X1_468/Y gnd OAI21X1_511/B vdd NAND2X1
XNAND2X1_453 AOI22X1_55/A AOI22X1_55/B gnd NAND3X1_506/B vdd NAND2X1
XNAND2X1_420 AOI22X1_49/A AOI22X1_49/B gnd NAND3X1_444/A vdd NAND2X1
XNAND2X1_464 OAI21X1_445/Y OR2X2_51/Y gnd XNOR2X1_50/B vdd NAND2X1
XNAND2X1_431 XOR2X1_33/Y INVX1_331/A gnd NAND3X1_495/B vdd NAND2X1
XNAND2X1_442 OR2X2_46/B OR2X2_46/A gnd NAND2X1_443/A vdd NAND2X1
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_52 NOR3X1_2/Y NOR2X1_48/B INVX1_78/Y gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_30 NOR2X1_40/A INVX1_58/Y INVX1_39/A gnd INVX1_59/A vdd OAI21X1
XOAI21X1_41 INVX1_16/Y INVX1_28/Y NOR2X1_46/A gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_63 INVX1_36/Y INVX1_18/Y OR2X2_13/A gnd OAI21X1_64/C vdd OAI21X1
XOAI21X1_74 NOR3X1_4/B NOR3X1_4/C OAI21X1_74/C gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_85 NOR3X1_12/B NOR3X1_12/C NOR3X1_12/A gnd OAI21X1_85/Y vdd OAI21X1
XOAI21X1_96 NOR2X1_46/B NOR2X1_76/A AOI22X1_9/A gnd OR2X2_15/A vdd OAI21X1
XOAI21X1_233 OAI21X1_234/A NOR3X1_21/Y INVX1_211/A gnd OAI21X1_233/Y vdd OAI21X1
XOAI21X1_255 OAI22X1_8/C INVX1_18/Y INVX1_195/Y gnd OAI21X1_256/C vdd OAI21X1
XOAI21X1_244 INVX1_185/Y NOR2X1_99/A INVX1_186/A gnd XOR2X1_15/B vdd OAI21X1
XOAI21X1_200 OAI21X1_200/A NOR3X1_20/Y INVX1_188/A gnd OAI21X1_200/Y vdd OAI21X1
XOAI21X1_222 OAI21X1_222/A AOI21X1_93/C INVX1_213/A gnd OAI21X1_237/C vdd OAI21X1
XOAI21X1_211 INVX1_168/Y XNOR2X1_30/B INVX1_170/Y gnd INVX1_196/A vdd OAI21X1
XAND2X2_99 OR2X2_47/A OR2X2_47/B gnd AND2X2_99/Y vdd AND2X2
XINVX1_308 INVX1_308/A gnd INVX1_308/Y vdd INVX1
XAND2X2_66 INVX1_261/Y AND2X2_66/B gnd INVX1_263/A vdd AND2X2
XAND2X2_77 AND2X2_77/A AND2X2_77/B gnd AND2X2_77/Y vdd AND2X2
XOAI21X1_288 NOR3X1_24/A NOR3X1_24/B OAI21X1_288/C gnd OAI21X1_288/Y vdd OAI21X1
XOAI21X1_277 INVX1_28/Y OAI22X1_6/D OAI21X1_277/C gnd OAI21X1_278/C vdd OAI21X1
XINVX1_319 vertices[13] gnd INVX1_319/Y vdd INVX1
XOAI21X1_299 NOR3X1_25/B NOR3X1_25/C NOR3X1_25/A gnd OAI21X1_299/Y vdd OAI21X1
XAND2X2_88 AND2X2_88/A AND2X2_88/B gnd XOR2X1_26/A vdd AND2X2
XAND2X2_44 INVX1_1/A vertices[9] gnd AND2X2_44/Y vdd AND2X2
XAND2X2_33 INVX1_109/A AND2X2_33/B gnd NOR3X1_6/A vdd AND2X2
XAND2X2_22 vertices[2] cos_alpha[4] gnd AND2X2_22/Y vdd AND2X2
XAND2X2_11 OR2X2_6/Y AOI21X1_1/B gnd XOR2X1_4/A vdd AND2X2
XAND2X2_55 OR2X2_25/Y AND2X2_59/A gnd AND2X2_55/Y vdd AND2X2
XOAI21X1_266 INVX1_202/A OAI21X1_266/B INVX1_248/A gnd OAI21X1_294/C vdd OAI21X1
XNAND2X1_283 OAI21X1_270/Y INVX1_242/Y gnd XOR2X1_18/B vdd NAND2X1
XNAND2X1_294 BUFX2_4/Y vertices[11] gnd NOR2X1_149/A vdd NAND2X1
XNAND2X1_250 AOI22X1_39/A AOI22X1_39/B gnd XOR2X1_16/A vdd NAND2X1
XNAND2X1_261 INVX1_233/Y OAI21X1_261/Y gnd AND2X2_67/B vdd NAND2X1
XNAND2X1_272 INVX1_236/A INVX1_237/A gnd NAND3X1_317/B vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XINVX1_116 NOR2X1_68/Y gnd OAI22X1_5/A vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XINVX1_138 NOR2X1_83/Y gnd OAI22X1_5/B vdd INVX1
XINVX1_149 NOR2X1_74/B gnd INVX1_149/Y vdd INVX1
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 NAND3X1_190/C NAND3X1_190/A OAI21X1_193/C gnd OAI21X1_220/B vdd AOI21X1
XFILL_18_2 gnd vdd FILL
XNAND3X1_66 INVX1_134/A INVX1_135/A NAND3X1_66/C gnd INVX1_111/A vdd NAND3X1
XNAND3X1_55 OAI21X1_76/Y INVX1_105/A OAI21X1_78/C gnd NAND3X1_59/C vdd NAND3X1
XNAND3X1_22 INVX1_77/A INVX1_104/A OAI21X1_50/Y gnd NAND3X1_22/Y vdd NAND3X1
XNAND3X1_33 NOR3X1_12/A AOI22X1_4/A INVX1_88/Y gnd INVX1_89/A vdd NAND3X1
XNAND3X1_11 INVX1_61/Y INVX1_60/A OAI21X1_33/Y gnd INVX1_88/A vdd NAND3X1
XNAND3X1_44 BUFX2_16/Y vertices[5] NOR2X1_58/B gnd NAND3X1_44/Y vdd NAND3X1
XNAND3X1_88 INVX1_98/A INVX1_156/A NAND3X1_88/C gnd NAND3X1_93/A vdd NAND3X1
XNOR2X1_66 NOR3X1_12/B NOR3X1_12/C gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_99 NOR2X1_99/A NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_11 OAI21X1_5/A XNOR2X1_1/Y gnd INVX1_14/A vdd NOR2X1
XNOR2X1_88 dy[8] dx[8] gnd NOR2X1_89/A vdd NOR2X1
XNAND3X1_77 NAND3X1_77/A NAND3X1_77/B NAND3X1_77/C gnd NAND3X1_81/B vdd NAND3X1
XNOR2X1_55 OR2X2_9/B OR2X2_9/A gnd NOR2X1_55/Y vdd NOR2X1
XNAND3X1_99 NOR2X1_73/A NAND3X1_99/B NAND3X1_99/C gnd NAND3X1_99/Y vdd NAND3X1
XNOR2X1_44 INVX1_41/Y INVX1_43/Y gnd INVX1_70/A vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_34/B vdd NOR2X1
XNOR2X1_22 NOR2X1_22/A INVX1_21/Y gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_77 NOR2X1_77/A NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XNAND3X1_499 INVX1_330/Y INVX1_385/A OAI21X1_470/Y gnd NAND3X1_502/A vdd NAND3X1
XNAND3X1_466 INVX1_354/Y NAND3X1_469/B NAND3X1_469/C gnd AOI22X1_53/C vdd NAND3X1
XNAND3X1_488 OAI21X1_463/Y OAI21X1_462/Y INVX1_341/Y gnd NAND3X1_492/A vdd NAND3X1
XNAND3X1_444 NAND3X1_444/A AOI22X1_48/C AOI22X1_48/D gnd AND2X2_102/A vdd NAND3X1
XNAND3X1_422 NAND3X1_424/A NAND3X1_425/B OAI21X1_405/Y gnd NAND3X1_423/C vdd NAND3X1
XNAND3X1_400 INVX1_307/A NAND3X1_436/B NAND3X1_436/C gnd AOI22X1_46/A vdd NAND3X1
XNAND3X1_411 OAI21X1_395/Y NAND3X1_411/B OAI21X1_396/Y gnd INVX1_320/A vdd NAND3X1
XNAND3X1_433 INVX1_308/A AOI22X1_45/C AOI22X1_45/D gnd NAND3X1_434/C vdd NAND3X1
XNAND3X1_477 AND2X2_79/Y INVX1_323/A AOI22X1_41/Y gnd NAND3X1_481/B vdd NAND3X1
XNAND3X1_455 INVX1_336/A INVX1_337/A INVX1_338/Y gnd NAND3X1_455/Y vdd NAND3X1
XNOR2X1_178 NOR2X1_178/A NOR2X1_178/B gnd NOR2X1_179/B vdd NOR2X1
XNOR2X1_189 INVX1_372/Y XNOR2X1_73/Y gnd OAI22X1_10/A vdd NOR2X1
XNOR2X1_145 OR2X2_33/B OR2X2_33/A gnd NOR3X1_26/C vdd NOR2X1
XNOR2X1_123 XOR2X1_19/B XOR2X1_19/A gnd OR2X2_34/A vdd NOR2X1
XNOR2X1_167 INVX1_334/Y XNOR2X1_40/A gnd OR2X2_45/A vdd NOR2X1
XNOR2X1_112 INVX1_91/Y OAI22X1_8/D gnd NOR2X1_113/B vdd NOR2X1
XNOR2X1_134 NOR2X1_134/A INVX1_266/Y gnd OR2X2_30/A vdd NOR2X1
XNOR2X1_156 NOR2X1_91/A OAI22X1_8/D gnd INVX1_334/A vdd NOR2X1
XNOR2X1_101 INVX1_91/Y OAI22X1_8/B gnd INVX1_229/A vdd NOR2X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_25 XOR2X1_1/Y gnd INVX1_25/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_36 cos_gamma[4] gnd INVX1_36/Y vdd INVX1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XNAND3X1_230 XNOR2X1_32/Y OAI21X1_233/Y OAI21X1_276/C gnd NAND3X1_235/A vdd NAND3X1
XNAND3X1_241 INVX1_247/A OAI21X1_238/Y INVX1_214/Y gnd NAND3X1_244/B vdd NAND3X1
XNAND3X1_285 NOR2X1_121/Y INVX1_281/A OAI21X1_328/C gnd NAND3X1_285/Y vdd NAND3X1
XNAND3X1_296 NAND3X1_298/A OAI21X1_290/Y OAI21X1_291/C gnd NAND3X1_297/C vdd NAND3X1
XNAND3X1_274 AOI22X1_38/A NAND3X1_276/A NAND3X1_276/B gnd INVX1_256/A vdd NAND3X1
XNAND3X1_252 INVX1_201/Y NAND3X1_252/B NAND3X1_252/C gnd NAND3X1_255/C vdd NAND3X1
XNAND3X1_263 INVX1_222/A INVX1_221/Y NAND3X1_263/C gnd NAND3X1_264/A vdd NAND3X1
XOAI21X1_437 INVX1_73/Y NOR2X1_95/B OAI21X1_437/C gnd OAI21X1_438/C vdd OAI21X1
XOAI21X1_404 OAI21X1_430/B NOR3X1_41/Y INVX1_322/Y gnd OAI21X1_404/Y vdd OAI21X1
XOAI21X1_415 AOI22X1_50/Y AOI22X1_51/Y OAI21X1_415/C gnd OAI21X1_415/Y vdd OAI21X1
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_448 INVX1_71/Y OAI22X1_6/B OR2X2_52/A gnd OAI21X1_448/Y vdd OAI21X1
XOAI21X1_426 OR2X2_37/A INVX1_342/Y OAI21X1_426/C gnd INVX1_346/A vdd OAI21X1
XOAI21X1_459 INVX1_324/Y NOR2X1_162/A INVX1_325/A gnd XOR2X1_39/B vdd OAI21X1
XNAND2X1_454 NAND3X1_405/B NAND3X1_405/Y gnd XNOR2X1_48/A vdd NAND2X1
XNAND2X1_487 AND2X2_96/B AND2X2_96/A gnd NAND3X1_505/A vdd NAND2X1
XNAND2X1_498 NAND3X1_510/A NAND3X1_510/B gnd NAND2X1_499/B vdd NAND2X1
XNAND2X1_476 XOR2X1_36/Y OAI21X1_483/B gnd NAND3X1_469/C vdd NAND2X1
XNAND2X1_432 INVX1_332/Y INVX1_331/Y gnd NAND3X1_495/C vdd NAND2X1
XNAND2X1_421 OR2X2_41/B OR2X2_41/A gnd AOI22X1_51/B vdd NAND2X1
XNAND2X1_443 NAND2X1_443/A OR2X2_46/Y gnd XNOR2X1_47/A vdd NAND2X1
XNAND2X1_410 INVX1_323/Y OAI21X1_406/Y gnd NAND2X1_411/B vdd NAND2X1
XNAND2X1_465 cos_alpha[4] vertices[11] gnd OR2X2_57/B vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XOAI21X1_53 NOR3X1_2/Y NOR2X1_48/B INVX1_78/A gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_42 NOR2X1_46/Y NOR2X1_47/Y INVX1_72/Y gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_86 INVX1_63/A NOR2X1_52/A INVX1_89/A gnd XNOR2X1_17/B vdd OAI21X1
XOAI21X1_75 OAI21X1_75/A OAI21X1_75/B OAI21X1_75/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_31 INVX1_59/Y AND2X2_14/Y INVX1_35/A gnd AOI21X1_6/A vdd OAI21X1
XOAI21X1_64 OAI21X1_64/A OAI21X1_91/C OAI21X1_64/C gnd XNOR2X1_15/A vdd OAI21X1
XOAI21X1_20 INVX1_36/Y INVX1_9/Y OAI21X1_36/A gnd OAI21X1_21/C vdd OAI21X1
XOAI21X1_97 OAI21X1_97/A OAI21X1_97/B AOI22X1_9/C gnd OAI21X1_97/Y vdd OAI21X1
XOAI21X1_223 INVX1_29/Y INVX1_146/Y NOR2X1_142/A gnd OAI21X1_224/C vdd OAI21X1
XOAI21X1_278 NOR2X1_146/A AND2X2_75/A OAI21X1_278/C gnd XOR2X1_20/A vdd OAI21X1
XOAI21X1_289 OAI21X1_291/A OAI21X1_291/B OAI21X1_289/C gnd OAI21X1_289/Y vdd OAI21X1
XOAI21X1_256 OAI21X1_311/A OAI21X1_314/C OAI21X1_256/C gnd INVX1_228/A vdd OAI21X1
XOAI21X1_234 OAI21X1_234/A NOR3X1_21/Y INVX1_211/Y gnd OAI21X1_234/Y vdd OAI21X1
XOAI21X1_267 INVX1_214/A OAI21X1_267/B INVX1_247/A gnd OAI21X1_293/C vdd OAI21X1
XOAI21X1_212 NOR2X1_91/A INVX1_18/Y INVX1_197/Y gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_201 AOI22X1_25/Y OAI21X1_202/B INVX1_189/A gnd OAI21X1_201/Y vdd OAI21X1
XOAI21X1_245 OAI21X1_246/A INVX1_222/Y INVX1_221/Y gnd AOI22X1_28/D vdd OAI21X1
XINVX1_309 INVX1_309/A gnd OR2X2_48/A vdd INVX1
XAND2X2_89 AND2X2_89/A AND2X2_89/B gnd AND2X2_89/Y vdd AND2X2
XAND2X2_67 AND2X2_67/A AND2X2_67/B gnd INVX1_262/A vdd AND2X2
XAND2X2_78 AND2X2_78/A INVX1_239/A gnd AND2X2_78/Y vdd AND2X2
XAND2X2_23 vertices[3] cos_alpha[3] gnd AND2X2_23/Y vdd AND2X2
XAND2X2_34 INVX1_139/Y AND2X2_34/B gnd INVX1_140/A vdd AND2X2
XAND2X2_12 BUFX2_15/Y vertices[4] gnd AOI22X1_2/B vdd AND2X2
XAND2X2_45 OR2X2_21/Y INVX1_202/A gnd AND2X2_45/Y vdd AND2X2
XAND2X2_56 AND2X2_56/A AND2X2_56/B gnd AND2X2_56/Y vdd AND2X2
XNAND2X1_295 NAND3X1_292/Y NAND3X1_293/Y gnd OAI21X1_331/B vdd NAND2X1
XNAND2X1_284 NAND3X1_233/A NAND3X1_233/Y gnd XOR2X1_18/A vdd NAND2X1
XNAND2X1_251 INVX1_255/A NAND3X1_276/A gnd OAI21X1_307/C vdd NAND2X1
XNAND2X1_262 INVX1_233/A AND2X2_61/Y gnd NAND3X1_324/C vdd NAND2X1
XNAND2X1_240 OAI21X1_242/C OAI21X1_354/A gnd NAND2X1_242/B vdd NAND2X1
XNAND2X1_273 INVX1_237/A INVX1_236/Y gnd NAND3X1_318/B vdd NAND2X1
XFILL_26_0_1 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XINVX1_106 dz[6] gnd INVX1_106/Y vdd INVX1
XINVX1_117 NOR2X1_69/Y gnd NOR3X1_17/A vdd INVX1
XINVX1_139 NOR2X1_84/Y gnd INVX1_139/Y vdd INVX1
XINVX1_128 vertices[7] gnd INVX1_128/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XNAND3X1_89 OR2X2_10/A NAND3X1_89/B NAND3X1_89/C gnd NAND3X1_93/C vdd NAND3X1
XNAND3X1_67 INVX1_113/Y INVX1_112/Y OR2X2_12/Y gnd NAND3X1_68/B vdd NAND3X1
XNOR2X1_12 INVX1_6/Y AND2X2_4/A gnd NOR2X1_13/A vdd NOR2X1
XNAND3X1_23 OAI21X1_47/Y INVX1_76/A OAI21X1_50/C gnd NAND3X1_37/C vdd NAND3X1
XNAND3X1_56 OAI21X1_79/Y NAND3X1_58/C NAND3X1_59/C gnd NAND3X1_57/B vdd NAND3X1
XNAND3X1_45 NOR3X1_4/A NAND3X1_45/B OAI21X1_72/Y gnd NAND3X1_46/B vdd NAND3X1
XNAND3X1_78 NAND3X1_78/A NAND3X1_78/B NAND3X1_78/C gnd NAND3X1_81/A vdd NAND3X1
XNAND3X1_34 INVX1_94/A NAND3X1_34/B OR2X2_9/Y gnd AND2X2_21/B vdd NAND3X1
XNAND3X1_12 NOR2X1_29/Y INVX1_88/A AOI21X1_8/A gnd INVX1_63/A vdd NAND3X1
XNAND3X1_423 NAND3X1_423/A INVX1_358/A NAND3X1_423/C gnd NAND3X1_423/Y vdd NAND3X1
XNAND3X1_401 INVX1_307/Y NAND3X1_437/B NAND3X1_437/C gnd AOI22X1_46/B vdd NAND3X1
XNAND3X1_412 OAI21X1_395/C NAND3X1_412/B NAND3X1_412/C gnd NAND3X1_413/C vdd NAND3X1
XNOR2X1_89 NOR2X1_89/A NOR2X1_89/B gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_56 INVX1_41/Y OAI22X1_8/B gnd INVX1_96/A vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd INVX1_38/A vdd NOR2X1
XNOR2X1_45 INVX1_2/Y INVX1_71/Y gnd INVX1_72/A vdd NOR2X1
XNOR2X1_23 NOR2X1_43/A INVX1_23/Y gnd INVX1_24/A vdd NOR2X1
XNOR2X1_78 NOR2X1_78/A NOR2X1_78/B gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_83/A NOR2X1_7/B gnd NOR2X1_67/Y vdd NOR2X1
XNAND3X1_467 AOI22X1_53/D AOI22X1_53/C AND2X2_101/Y gnd NAND3X1_473/C vdd NAND3X1
XNAND3X1_445 OAI21X1_414/C NAND3X1_446/A AND2X2_102/A gnd AOI22X1_50/C vdd NAND3X1
XNAND3X1_456 INVX1_339/Y NAND3X1_456/B OR2X2_47/Y gnd NAND3X1_456/Y vdd NAND3X1
XNAND3X1_489 INVX1_341/A OAI21X1_464/Y OAI21X1_465/Y gnd NAND3X1_492/B vdd NAND3X1
XNAND3X1_434 XOR2X1_31/Y NAND3X1_434/B NAND3X1_434/C gnd AOI22X1_55/B vdd NAND3X1
XNAND3X1_478 OAI21X1_458/C NAND3X1_481/B NAND3X1_478/C gnd NAND3X1_478/Y vdd NAND3X1
XNOR2X1_102 NOR2X1_102/A NOR2X1_140/A gnd INVX1_204/A vdd NOR2X1
XNOR2X1_124 INVX1_71/Y INVX1_177/Y gnd XOR2X1_20/B vdd NOR2X1
XNOR2X1_113 NOR2X1_113/A NOR2X1_113/B gnd NOR2X1_115/B vdd NOR2X1
XNOR2X1_179 NOR2X1_179/A NOR2X1_179/B gnd NOR2X1_179/Y vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XNOR2X1_135 AND2X2_71/B AND2X2_71/A gnd NOR2X1_136/A vdd NOR2X1
XNOR2X1_146 NOR2X1_146/A AND2X2_75/A gnd NOR2X1_146/Y vdd NOR2X1
XNOR2X1_157 INVX1_22/Y NOR2X1_197/B gnd NOR2X1_157/Y vdd NOR2X1
XNOR2X1_168 NOR2X1_91/A INVX1_124/Y gnd INVX1_336/A vdd NOR2X1
XINVX1_26 INVX1_26/A gnd OR2X2_6/B vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XAOI21X1_260 OAI21X1_507/Y NAND3X1_536/B XNOR2X1_59/Y gnd NOR3X1_50/A vdd AOI21X1
XNAND3X1_231 OAI21X1_236/C NAND3X1_235/A OAI21X1_232/Y gnd INVX1_246/A vdd NAND3X1
XNAND3X1_220 NOR3X1_19/C NAND3X1_275/A OAI21X1_205/Y gnd OAI21X1_308/C vdd NAND3X1
XNAND3X1_275 NAND3X1_275/A INVX1_256/A OAI21X1_251/Y gnd AOI22X1_39/A vdd NAND3X1
XNAND3X1_264 NAND3X1_264/A NAND3X1_264/B OAI21X1_246/Y gnd NAND3X1_268/B vdd NAND3X1
XNAND3X1_253 INVX1_216/Y NAND3X1_255/B NAND3X1_255/C gnd AOI22X1_32/B vdd NAND3X1
XNAND3X1_242 INVX1_215/A NAND3X1_244/A NAND3X1_244/B gnd INVX1_248/A vdd NAND3X1
XNAND3X1_286 OR2X2_29/Y OAI21X1_275/Y NAND3X1_293/C gnd NAND3X1_286/Y vdd NAND3X1
XNAND3X1_297 XOR2X1_18/Y OAI21X1_289/Y NAND3X1_297/C gnd NAND3X1_301/A vdd NAND3X1
XOAI21X1_438 OAI21X1_486/A XNOR2X1_64/A OAI21X1_438/C gnd OR2X2_49/A vdd OAI21X1
XOAI21X1_405 OAI21X1_430/B NOR3X1_41/Y INVX1_322/A gnd OAI21X1_405/Y vdd OAI21X1
XOAI21X1_416 AOI22X1_50/Y AOI22X1_51/Y AND2X2_94/Y gnd AOI22X1_52/D vdd OAI21X1
XFILL_21_1_2 gnd vdd FILL
XOAI21X1_449 AND2X2_90/Y INVX1_318/Y OR2X2_40/Y gnd XOR2X1_37/B vdd OAI21X1
XOAI21X1_427 INVX1_343/A INVX1_345/Y INVX1_344/Y gnd AND2X2_100/A vdd OAI21X1
XNAND2X1_400 INVX1_316/Y OAI21X1_440/A gnd NAND3X1_408/C vdd NAND2X1
XNAND2X1_411 NAND3X1_427/Y NAND2X1_411/B gnd NAND3X1_432/C vdd NAND2X1
XNAND2X1_455 vertices[2] cos_alpha[13] gnd XNOR2X1_63/A vdd NAND2X1
XNAND2X1_477 AOI22X1_53/A AOI22X1_53/B gnd OAI21X1_497/B vdd NAND2X1
XNAND2X1_488 AOI22X1_56/B AOI22X1_56/A gnd NOR2X1_178/A vdd NAND2X1
XNAND2X1_499 XNOR2X1_61/Y NAND2X1_499/B gnd NAND3X1_533/A vdd NAND2X1
XNAND2X1_444 OR2X2_47/B OR2X2_47/A gnd NAND3X1_456/B vdd NAND2X1
XNAND2X1_422 AOI22X1_51/B OR2X2_41/Y gnd INVX1_328/A vdd NAND2X1
XNAND2X1_433 NAND3X1_495/B NAND3X1_495/C gnd XNOR2X1_46/A vdd NAND2X1
XNAND2X1_466 cos_alpha[5] vertices[9] gnd OR2X2_52/B vdd NAND2X1
XFILL_4_2_2 gnd vdd FILL
XFILL_12_1_2 gnd vdd FILL
XOAI21X1_87 INVX1_93/A NOR2X1_64/A INVX1_111/A gnd OAI21X1_87/Y vdd OAI21X1
XOAI21X1_10 NOR2X1_9/A NOR2X1_9/B AND2X2_2/B gnd OR2X2_4/A vdd OAI21X1
XOAI21X1_76 OAI21X1_95/B NOR3X1_3/Y OR2X2_10/Y gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_54 INVX1_79/A OAI21X1_54/B INVX1_70/Y gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_65 NOR2X1_55/Y AND2X2_20/Y INVX1_94/Y gnd AND2X2_21/A vdd OAI21X1
XOAI21X1_32 NOR2X1_42/A INVX1_60/Y INVX1_61/A gnd AOI21X1_8/A vdd OAI21X1
XOAI21X1_98 INVX1_28/Y INVX1_50/Y NOR2X1_76/A gnd OAI21X1_98/Y vdd OAI21X1
XOAI21X1_21 NOR2X1_43/A INVX1_37/Y OAI21X1_21/C gnd NOR2X1_34/A vdd OAI21X1
XOAI21X1_43 INVX1_1/Y INVX1_73/Y OAI21X1_43/C gnd AOI22X1_7/D vdd OAI21X1
XOAI21X1_268 INVX1_45/Y INVX1_203/Y OAI21X1_325/A gnd OAI21X1_269/C vdd OAI21X1
XOAI21X1_257 INVX1_226/Y INVX1_9/Y INVX1_228/A gnd AND2X2_60/B vdd OAI21X1
XOAI21X1_224 OAI21X1_224/A OAI21X1_272/C OAI21X1_224/C gnd XOR2X1_13/A vdd OAI21X1
XOAI21X1_279 NOR3X1_21/A NOR3X1_21/C OAI21X1_279/C gnd OAI21X1_286/C vdd OAI21X1
XOAI21X1_235 OAI21X1_236/A OAI21X1_236/B OAI21X1_235/C gnd OAI21X1_235/Y vdd OAI21X1
XAND2X2_13 NAND3X1_8/Y NOR2X1_60/A gnd AND2X2_13/Y vdd AND2X2
XOAI21X1_202 AOI22X1_25/Y OAI21X1_202/B INVX1_189/Y gnd AOI22X1_26/D vdd OAI21X1
XOAI21X1_213 INVX1_172/Y NOR2X1_94/Y OAI21X1_213/C gnd XNOR2X1_31/A vdd OAI21X1
XOAI21X1_246 OAI21X1_246/A INVX1_222/Y INVX1_221/A gnd OAI21X1_246/Y vdd OAI21X1
XAND2X2_79 AND2X2_79/A INVX1_359/A gnd AND2X2_79/Y vdd AND2X2
XAND2X2_68 AND2X2_82/B AND2X2_68/B gnd INVX1_265/A vdd AND2X2
XNAND2X1_230 cos_alpha[3] vertices[6] gnd OAI21X1_229/A vdd NAND2X1
XAND2X2_35 OR2X2_16/Y AND2X2_35/B gnd AND2X2_35/Y vdd AND2X2
XAND2X2_57 INVX1_192/A AND2X2_57/B gnd AND2X2_57/Y vdd AND2X2
XAND2X2_24 BUFX2_15/Y vertices[6] gnd AND2X2_24/Y vdd AND2X2
XAND2X2_46 AND2X2_46/A AND2X2_46/B gnd AND2X2_46/Y vdd AND2X2
XNAND2X1_252 XNOR2X1_31/A AND2X2_58/Y gnd AND2X2_59/B vdd NAND2X1
XNAND2X1_241 INVX1_239/A NAND3X1_255/Y gnd OAI21X1_354/B vdd NAND2X1
XNAND2X1_285 vertices[3] cos_alpha[8] gnd XOR2X1_19/B vdd NAND2X1
XNAND2X1_296 AND2X2_78/A AND2X2_64/A gnd OAI21X1_296/C vdd NAND2X1
XNAND2X1_263 INVX1_233/Y AND2X2_61/Y gnd NAND3X1_325/C vdd NAND2X1
XNAND2X1_274 INVX1_236/A INVX1_237/Y gnd NAND3X1_318/C vdd NAND2X1
XFILL_26_0_2 gnd vdd FILL
XFILL_1_0_2 gnd vdd FILL
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_107 INVX1_107/A gnd NOR2X1_63/B vdd INVX1
XINVX1_129 OR2X2_11/A gnd INVX1_129/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XFILL_17_0_2 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XNAND3X1_35 cos_gamma[1] OAI21X1_53/Y NAND3X1_35/C gnd OR2X2_11/B vdd NAND3X1
XNAND3X1_57 NAND3X1_57/A NAND3X1_57/B NAND3X1_57/C gnd NAND3X1_61/B vdd NAND3X1
XNAND3X1_79 NAND3X1_81/B NAND3X1_81/A NOR3X1_14/C gnd NAND3X1_80/B vdd NAND3X1
XNAND3X1_68 OAI21X1_85/Y NAND3X1_68/B XNOR2X1_17/B gnd XNOR2X1_19/B vdd NAND3X1
XNOR2X1_13 NOR2X1_13/A AND2X2_4/Y gnd NOR2X1_13/Y vdd NOR2X1
XNAND3X1_46 OAI21X1_97/A NAND3X1_46/B OAI21X1_74/Y gnd NAND3X1_50/A vdd NAND3X1
XNAND3X1_24 INVX1_77/Y OAI21X1_51/Y NAND3X1_37/C gnd NAND3X1_24/Y vdd NAND3X1
XNOR2X1_46 NOR2X1_46/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_35 INVX1_41/Y INVX1_18/Y gnd INVX1_42/A vdd NOR2X1
XNOR2X1_24 AND2X2_8/B AND2X2_8/A gnd NOR2X1_25/A vdd NOR2X1
XNAND3X1_13 cos_gamma[5] INVX1_9/A INVX1_66/Y gnd OAI21X1_62/C vdd NAND3X1
XNAND3X1_402 INVX1_311/Y NAND3X1_402/B NAND3X1_402/C gnd OAI21X1_432/C vdd NAND3X1
XNAND3X1_446 NAND3X1_446/A AND2X2_102/A AND2X2_93/Y gnd AOI22X1_51/C vdd NAND3X1
XNAND3X1_435 INVX1_327/A AOI22X1_55/B OAI21X1_408/Y gnd INVX1_340/A vdd NAND3X1
XNAND3X1_424 NAND3X1_424/A NAND3X1_424/B OAI21X1_404/Y gnd NAND3X1_426/B vdd NAND3X1
XNAND3X1_413 XNOR2X1_44/Y INVX1_320/A NAND3X1_413/C gnd NAND3X1_414/B vdd NAND3X1
XNAND3X1_457 cos_gamma[5] NAND3X1_457/B XOR2X1_26/A gnd OAI21X1_426/C vdd NAND3X1
XNOR2X1_57 INVX1_97/Y NOR2X1_57/B gnd OR2X2_10/B vdd NOR2X1
XNOR2X1_79 dy[7] dx[7] gnd NOR2X1_80/A vdd NOR2X1
XNOR2X1_68 INVX1_91/Y NOR2X1_7/B gnd NOR2X1_68/Y vdd NOR2X1
XNAND3X1_468 INVX1_354/Y NAND3X1_468/B NAND3X1_468/C gnd NAND3X1_470/A vdd NAND3X1
XNAND3X1_479 AND2X2_79/A INVX1_359/A INVX1_323/A gnd OAI21X1_458/B vdd NAND3X1
XNOR2X1_158 XOR2X1_23/A XOR2X1_23/B gnd NOR2X1_158/Y vdd NOR2X1
XNOR2X1_136 NOR2X1_136/A AND2X2_71/Y gnd NOR2X1_136/Y vdd NOR2X1
XNOR2X1_114 INVX1_229/Y NOR2X1_133/A gnd NOR2X1_115/A vdd NOR2X1
XNOR2X1_103 XOR2X1_13/B XOR2X1_13/A gnd OR2X2_29/A vdd NOR2X1
XNOR2X1_125 AND2X2_51/B NOR2X1_125/B gnd NOR2X1_125/Y vdd NOR2X1
XNOR2X1_147 INVX1_71/Y INVX1_128/Y gnd INVX1_285/A vdd NOR2X1
XFILL_23_2 gnd vdd FILL
XFILL_16_1 gnd vdd FILL
XNOR2X1_169 NOR2X1_169/A XNOR2X1_79/A gnd INVX1_338/A vdd NOR2X1
XINVX1_27 NOR2X1_7/B gnd INVX1_27/Y vdd INVX1
XINVX1_290 NOR3X1_34/A gnd INVX1_290/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XINVX1_16 vertices[2] gnd INVX1_16/Y vdd INVX1
XFILL_24_1_0 gnd vdd FILL
XNAND2X1_90 BUFX2_4/Y vertices[6] gnd NOR2X1_58/B vdd NAND2X1
XAOI21X1_250 NAND3X1_521/C NAND3X1_521/B NAND3X1_523/A gnd OAI22X1_13/A vdd AOI21X1
XAOI21X1_261 AOI22X1_59/D AOI22X1_59/C INVX1_382/Y gnd NOR3X1_51/B vdd AOI21X1
XFILL_7_2_0 gnd vdd FILL
XNAND3X1_287 INVX1_244/Y OAI21X1_281/Y OAI21X1_340/C gnd NAND3X1_291/B vdd NAND3X1
XNAND3X1_298 NAND3X1_298/A OAI21X1_290/Y OAI21X1_289/C gnd INVX1_289/A vdd NAND3X1
XFILL_15_1_0 gnd vdd FILL
XNAND3X1_232 NAND3X1_232/A INVX1_211/A OAI21X1_230/Y gnd NAND3X1_232/Y vdd NAND3X1
XNAND3X1_210 INVX1_188/Y NAND3X1_210/B OAI21X1_198/Y gnd NAND3X1_211/B vdd NAND3X1
XNAND3X1_276 NAND3X1_276/A NAND3X1_276/B AND2X2_57/Y gnd NAND3X1_277/B vdd NAND3X1
XNAND3X1_254 INVX1_216/Y AOI22X1_41/A NAND3X1_254/C gnd INVX1_239/A vdd NAND3X1
XNAND3X1_243 INVX1_202/Y INVX1_248/A OAI21X1_239/Y gnd NAND3X1_251/B vdd NAND3X1
XNAND3X1_265 INVX1_253/A AOI22X1_28/D AND2X2_54/Y gnd NAND3X1_268/C vdd NAND3X1
XNAND3X1_221 OAI22X1_5/Y OAI21X1_168/Y INVX1_170/Y gnd NAND3X1_221/Y vdd NAND3X1
XOAI21X1_439 INVX1_29/Y INVX1_241/Y OR2X2_49/A gnd OAI21X1_439/Y vdd OAI21X1
XOAI21X1_417 NOR3X1_43/B NOR3X1_43/C NOR3X1_43/A gnd OAI21X1_417/Y vdd OAI21X1
XOAI21X1_428 NOR2X1_173/Y NOR3X1_42/C OAI21X1_428/C gnd OAI21X1_428/Y vdd OAI21X1
XOAI21X1_406 OAI21X1_406/A OAI21X1_458/A INVX1_359/A gnd OAI21X1_406/Y vdd OAI21X1
XNAND2X1_423 OAI21X1_472/C OAI21X1_417/Y gnd XOR2X1_32/A vdd NAND2X1
XNAND2X1_434 AOI22X1_48/C AND2X2_102/A gnd NAND3X1_498/A vdd NAND2X1
XNAND2X1_445 NAND3X1_456/Y OAI21X1_425/Y gnd INVX1_363/A vdd NAND2X1
XNAND2X1_401 INVX1_316/Y XOR2X1_28/Y gnd NAND3X1_409/B vdd NAND2X1
XNAND2X1_412 INVX1_323/A OAI21X1_406/Y gnd NAND3X1_508/C vdd NAND2X1
XNAND2X1_456 OAI21X1_435/Y OAI21X1_491/C gnd XOR2X1_35/B vdd NAND2X1
XNAND2X1_489 INVX1_385/A NAND3X1_502/A gnd OAI21X1_515/C vdd NAND2X1
XNAND2X1_478 OAI21X1_454/Y OAI21X1_455/Y gnd NAND3X1_478/C vdd NAND2X1
XNAND2X1_467 OAI21X1_448/Y OR2X2_52/Y gnd XNOR2X1_52/B vdd NAND2X1
XOAI21X1_11 XOR2X1_1/B XOR2X1_1/A NAND3X1_2/Y gnd INVX1_23/A vdd OAI21X1
XOAI21X1_66 INVX1_82/Y OAI21X1_66/B AND2X2_26/B gnd OAI21X1_66/Y vdd OAI21X1
XOAI21X1_77 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_55 INVX1_8/Y OAI22X1_8/B NOR2X1_49/B gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_22 OR2X2_5/B OR2X2_5/A OAI21X1_22/C gnd INVX1_40/A vdd OAI21X1
XOAI21X1_33 AOI21X1_7/Y INVX1_62/Y INVX1_24/Y gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_99 NOR2X1_76/Y NOR2X1_77/Y INVX1_126/A gnd OAI21X1_99/Y vdd OAI21X1
XOAI21X1_44 INVX1_10/Y INVX1_50/Y AND2X2_17/Y gnd OAI21X1_44/Y vdd OAI21X1
XOAI21X1_88 NOR2X1_83/A INVX1_9/Y OAI22X1_5/A gnd OAI21X1_89/C vdd OAI21X1
XOAI21X1_203 AOI22X1_26/Y OAI21X1_203/B INVX1_190/Y gnd OAI21X1_203/Y vdd OAI21X1
XOAI21X1_269 NOR2X1_140/A XOR2X1_23/A OAI21X1_269/C gnd XOR2X1_17/A vdd OAI21X1
XOAI21X1_225 OR2X2_29/A AND2X2_50/Y INVX1_206/Y gnd OAI21X1_225/Y vdd OAI21X1
XOAI21X1_258 XNOR2X1_30/B INVX1_229/Y OAI21X1_258/C gnd OAI21X1_258/Y vdd OAI21X1
XOAI21X1_236 OAI21X1_236/A OAI21X1_236/B OAI21X1_236/C gnd OAI21X1_236/Y vdd OAI21X1
XAND2X2_25 OR2X2_11/A OR2X2_11/B gnd AND2X2_25/Y vdd AND2X2
XAND2X2_14 NOR2X1_40/Y INVX1_39/Y gnd AND2X2_14/Y vdd AND2X2
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XAND2X2_47 OR2X2_17/Y AND2X2_47/B gnd AND2X2_47/Y vdd AND2X2
XOAI21X1_247 AOI22X1_28/Y OAI21X1_248/B OAI21X1_247/C gnd OAI21X1_247/Y vdd OAI21X1
XOAI21X1_214 OR2X2_19/B OR2X2_19/A AND2X2_40/B gnd INVX1_200/A vdd OAI21X1
XNAND2X1_220 vertices[0] cos_alpha[10] gnd NOR2X1_102/A vdd NAND2X1
XNAND2X1_286 vertices[5] cos_alpha[7] gnd OR2X2_32/A vdd NAND2X1
XAND2X2_69 AND2X2_69/A AND2X2_82/A gnd INVX1_267/A vdd AND2X2
XNAND2X1_231 cos_alpha[4] vertices[7] gnd OAI21X1_277/C vdd NAND2X1
XNAND2X1_253 INVX1_193/Y INVX1_195/A gnd OR2X2_27/B vdd NAND2X1
XNAND2X1_275 XOR2X1_15/B XOR2X1_15/A gnd AND2X2_65/B vdd NAND2X1
XAND2X2_58 OR2X2_24/Y AND2X2_58/B gnd AND2X2_58/Y vdd AND2X2
XNAND2X1_242 OAI21X1_241/Y NAND2X1_242/B gnd NAND3X1_256/C vdd NAND2X1
XNAND2X1_264 INVX1_233/A OAI21X1_261/Y gnd NAND3X1_325/B vdd NAND2X1
XNAND2X1_297 OAI21X1_296/Y NAND3X1_308/Y gnd AOI22X1_45/B vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNAND3X1_14 NOR2X1_43/Y NAND3X1_14/B OR2X2_8/Y gnd AND2X2_19/A vdd NAND3X1
XNAND3X1_25 BUFX2_5/Y OAI21X1_53/Y NAND3X1_35/C gnd NOR2X1_49/B vdd NAND3X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_47/B gnd NOR2X1_47/Y vdd NOR2X1
XNAND3X1_36 INVX1_77/Y INVX1_104/A OAI21X1_50/Y gnd NAND3X1_38/B vdd NAND3X1
XNAND3X1_58 INVX1_125/A OAI21X1_78/Y NAND3X1_58/C gnd NAND3X1_96/A vdd NAND3X1
XNOR2X1_14 INVX1_3/A INVX1_11/Y gnd XOR2X1_3/B vdd NOR2X1
XNAND3X1_69 INVX1_119/A INVX1_121/A INVX1_122/Y gnd AND2X2_27/A vdd NAND3X1
XNAND3X1_47 INVX1_99/A OAI22X1_4/Y NAND3X1_47/C gnd NAND3X1_47/Y vdd NAND3X1
XNOR2X1_25 NOR2X1_25/A AND2X2_8/Y gnd AND2X2_9/A vdd NOR2X1
XNOR2X1_69 NOR2X1_69/A NOR2X1_69/B gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_58 NOR2X1_58/A NOR2X1_58/B gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_36 OAI21X1_7/B INVX1_52/A gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_403 INVX1_311/A NAND3X1_403/B NAND3X1_403/C gnd NAND3X1_406/B vdd NAND3X1
XNAND3X1_469 INVX1_354/A NAND3X1_469/B NAND3X1_469/C gnd NAND3X1_470/B vdd NAND3X1
XNAND3X1_447 INVX1_328/Y AOI22X1_51/C AOI22X1_51/D gnd NAND3X1_451/B vdd NAND3X1
XNAND3X1_425 OAI21X1_379/Y NAND3X1_425/B OAI21X1_405/Y gnd NAND3X1_426/C vdd NAND3X1
XNAND3X1_414 OAI21X1_398/Y NAND3X1_414/B INVX1_321/Y gnd OAI21X1_441/C vdd NAND3X1
XNAND3X1_436 INVX1_307/Y NAND3X1_436/B NAND3X1_436/C gnd AOI22X1_47/A vdd NAND3X1
XNAND3X1_458 INVX1_344/A INVX1_345/A INVX1_343/Y gnd AND2X2_100/B vdd NAND3X1
XNOR2X1_148 AND2X2_75/A AND2X2_75/B gnd INVX1_286/A vdd NOR2X1
XNOR2X1_159 INVX1_15/Y OAI22X1_9/B gnd INVX1_318/A vdd NOR2X1
XNOR2X1_115 NOR2X1_115/A NOR2X1_115/B gnd NOR2X1_115/Y vdd NOR2X1
XNOR2X1_137 NOR2X1_137/A NOR2X1_137/B gnd NOR2X1_137/Y vdd NOR2X1
XNOR2X1_104 INVX1_73/Y INVX1_71/Y gnd XOR2X1_14/B vdd NOR2X1
XNOR2X1_126 AND2X2_52/Y AND2X2_63/Y gnd NOR2X1_126/Y vdd NOR2X1
XFILL_23_3 gnd vdd FILL
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XNAND2X1_80 cos_gamma[4] INVX1_43/A gnd OAI21X1_91/C vdd NAND2X1
XNAND2X1_91 AND2X2_17/Y AND2X2_24/Y gnd AOI22X1_8/D vdd NAND2X1
XINVX1_28 cos_alpha[3] gnd INVX1_28/Y vdd INVX1
XFILL_24_1_1 gnd vdd FILL
XAOI21X1_251 NAND3X1_523/C NAND3X1_523/B OAI21X1_482/Y gnd OAI22X1_13/B vdd AOI21X1
XAOI21X1_240 NAND3X1_505/B NAND3X1_505/C AND2X2_96/Y gnd INVX1_386/A vdd AOI21X1
XAOI21X1_262 OAI21X1_512/Y NAND3X1_541/B NOR2X1_200/A gnd OAI21X1_514/A vdd AOI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XNAND3X1_299 XNOR2X1_35/Y INVX1_289/A OAI21X1_291/Y gnd NAND3X1_301/B vdd NAND3X1
XNAND3X1_288 NAND3X1_291/B OAI21X1_286/C OAI21X1_280/Y gnd OAI21X1_337/C vdd NAND3X1
XNAND3X1_233 NAND3X1_233/A INVX1_207/Y OAI21X1_225/Y gnd NAND3X1_233/Y vdd NAND3X1
XNAND3X1_222 cos_gamma[8] INVX1_18/A INVX1_197/A gnd OAI21X1_258/C vdd NAND3X1
XNAND3X1_200 NAND3X1_200/A NAND3X1_200/B INVX1_216/A gnd NAND3X1_200/Y vdd NAND3X1
XNAND3X1_211 NAND3X1_211/A NAND3X1_211/B OAI21X1_200/Y gnd NAND3X1_215/B vdd NAND3X1
XNAND3X1_277 NOR3X1_22/Y NAND3X1_277/B OAI21X1_252/Y gnd AOI22X1_39/B vdd NAND3X1
XNAND3X1_266 NAND3X1_268/B AND2X2_53/Y NAND3X1_268/C gnd NAND3X1_267/B vdd NAND3X1
XNAND3X1_255 INVX1_216/A NAND3X1_255/B NAND3X1_255/C gnd NAND3X1_255/Y vdd NAND3X1
XNAND3X1_244 NAND3X1_244/A NAND3X1_244/B INVX1_215/Y gnd NAND3X1_248/B vdd NAND3X1
XOAI21X1_407 INVX1_292/Y NOR2X1_151/A INVX1_293/A gnd XOR2X1_31/B vdd OAI21X1
XOAI21X1_418 INVX1_303/A OAI21X1_418/B OAI21X1_418/C gnd INVX1_331/A vdd OAI21X1
XOAI21X1_429 NOR2X1_173/Y NOR3X1_42/C AND2X2_100/Y gnd OAI21X1_429/Y vdd OAI21X1
XNAND2X1_424 AOI22X1_50/C AND2X2_103/A gnd OAI21X1_471/C vdd NAND2X1
XNAND2X1_457 vertices[5] cos_alpha[10] gnd XNOR2X1_64/A vdd NAND2X1
XNAND2X1_413 NAND3X1_432/B NOR2X1_173/B gnd NAND3X1_431/C vdd NAND2X1
XNAND2X1_402 INVX1_316/A OAI21X1_440/A gnd NAND3X1_409/C vdd NAND2X1
XNAND2X1_435 XNOR2X1_41/B XNOR2X1_41/A gnd OAI21X1_421/C vdd NAND2X1
XNAND2X1_446 cos_gamma[5] NAND3X1_399/B gnd INVX1_344/A vdd NAND2X1
XNAND2X1_468 BUFX2_13/Y vertices[12] gnd OR2X2_56/B vdd NAND2X1
XNAND2X1_479 INVX1_377/A OAI21X1_457/Y gnd NAND3X1_481/C vdd NAND2X1
XOAI21X1_34 INVX1_24/Y AOI21X1_7/Y INVX1_62/A gnd INVX1_87/A vdd OAI21X1
XOAI21X1_23 NOR2X1_46/A INVX1_30/Y OAI22X1_2/Y gnd INVX1_47/A vdd OAI21X1
XOAI21X1_12 INVX1_22/Y INVX1_9/Y INVX1_23/Y gnd AND2X2_6/B vdd OAI21X1
XOAI21X1_45 INVX1_1/Y INVX1_73/Y AOI22X1_2/B gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_56 INVX1_55/Y NOR2X1_38/A INVX1_56/A gnd XOR2X1_6/B vdd OAI21X1
XOAI21X1_67 INVX1_77/A OAI21X1_67/B INVX1_104/A gnd OAI21X1_79/C vdd OAI21X1
XOAI21X1_78 OAI21X1_79/A INVX1_105/Y OAI21X1_78/C gnd OAI21X1_78/Y vdd OAI21X1
XOAI21X1_89 NOR2X1_82/A NOR2X1_82/B OAI21X1_89/C gnd NOR2X1_69/A vdd OAI21X1
XOAI21X1_226 OR2X2_29/A AND2X2_50/Y OAI22X1_7/Y gnd OAI21X1_226/Y vdd OAI21X1
XOAI21X1_237 OAI21X1_238/A OAI21X1_238/B OAI21X1_237/C gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_204 NOR2X1_84/A NOR2X1_84/B OAI21X1_207/B gnd OAI21X1_204/Y vdd OAI21X1
XOAI21X1_215 INVX1_36/Y INVX1_124/Y OAI21X1_263/A gnd OAI21X1_216/C vdd OAI21X1
XOAI21X1_259 NOR2X1_115/A NOR2X1_115/B INVX1_230/Y gnd OAI21X1_259/Y vdd OAI21X1
XAND2X2_26 AND2X2_26/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XAND2X2_15 vertices[1] cos_alpha[4] gnd NOR2X1_47/A vdd AND2X2
XAND2X2_48 AND2X2_48/A AND2X2_48/B gnd AND2X2_48/Y vdd AND2X2
XOAI21X1_248 AOI22X1_28/Y OAI21X1_248/B AND2X2_53/Y gnd AOI22X1_29/D vdd OAI21X1
XAND2X2_59 AND2X2_59/A AND2X2_59/B gnd OR2X2_27/A vdd AND2X2
XAND2X2_37 BUFX2_15/Y vertices[7] gnd NOR2X1_97/A vdd AND2X2
XNAND2X1_287 INVX1_243/Y XOR2X1_19/Y gnd OAI21X1_328/C vdd NAND2X1
XNAND2X1_232 cos_alpha[3] vertices[7] gnd NOR2X1_146/A vdd NAND2X1
XNAND2X1_276 cos_gamma[2] NAND3X1_399/B gnd INVX1_249/A vdd NAND2X1
XNAND2X1_298 AOI22X1_31/B NOR2X1_137/B gnd NAND3X1_312/B vdd NAND2X1
XNAND2X1_265 AND2X2_67/A AOI22X1_35/B gnd NAND3X1_323/B vdd NAND2X1
XNAND2X1_254 AOI22X1_37/A OR2X2_27/Y gnd INVX1_225/A vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_210 OAI21X1_217/Y OAI21X1_262/C gnd INVX1_199/A vdd NAND2X1
XNAND2X1_221 NAND3X1_183/B NAND3X1_183/Y gnd OR2X2_26/A vdd NAND2X1
XNAND2X1_243 OAI21X1_354/B OAI21X1_354/A gnd NAND3X1_257/C vdd NAND2X1
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XFILL_10_2_2 gnd vdd FILL
XNAND3X1_37 INVX1_77/A OAI21X1_51/Y NAND3X1_37/C gnd NAND3X1_38/C vdd NAND3X1
XNAND3X1_48 INVX1_99/Y OAI21X1_69/Y OAI21X1_70/Y gnd NAND3X1_48/Y vdd NAND3X1
XNAND3X1_15 INVX1_72/A OAI21X1_41/Y OAI21X1_68/C gnd NAND3X1_15/Y vdd NAND3X1
XNAND3X1_26 INVX1_70/A OAI21X1_55/Y INVX1_79/Y gnd NAND3X1_27/C vdd NAND3X1
XNOR2X1_48 NOR3X1_2/Y NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_37 dy[4] dx[4] gnd NOR2X1_38/A vdd NOR2X1
XNOR2X1_59 OR2X2_10/B OR2X2_10/A gnd NOR2X1_59/Y vdd NOR2X1
XNAND3X1_59 NAND3X1_59/A OAI21X1_79/Y NAND3X1_59/C gnd NAND3X1_60/B vdd NAND3X1
XNOR2X1_26 INVX1_2/Y INVX1_28/Y gnd INVX1_30/A vdd NOR2X1
XNOR2X1_15 OR2X2_3/A INVX1_9/Y gnd NOR2X1_17/A vdd NOR2X1
XNAND3X1_404 INVX1_313/A NAND3X1_406/B OAI21X1_432/C gnd NAND3X1_405/B vdd NAND3X1
XNAND3X1_448 INVX1_328/A AOI22X1_50/C AOI22X1_50/D gnd AND2X2_103/A vdd NAND3X1
XNAND3X1_415 OAI21X1_441/C OAI21X1_400/Y AND2X2_91/Y gnd NAND3X1_416/B vdd NAND3X1
XNAND3X1_426 NOR3X1_34/Y NAND3X1_426/B NAND3X1_426/C gnd NAND3X1_426/Y vdd NAND3X1
XNAND3X1_437 INVX1_307/A NAND3X1_437/B NAND3X1_437/C gnd AOI22X1_47/B vdd NAND3X1
XNAND3X1_459 INVX1_346/A NAND3X1_459/B OAI21X1_428/Y gnd OAI21X1_478/C vdd NAND3X1
XNOR2X1_127 dy[11] dx[11] gnd NOR2X1_128/A vdd NOR2X1
XNOR2X1_116 NOR2X1_116/A INVX1_231/Y gnd NOR2X1_116/Y vdd NOR2X1
XNOR2X1_138 INVX1_41/Y NOR2X1_197/B gnd INVX1_273/A vdd NOR2X1
XNOR2X1_149 NOR2X1_149/A OR2X2_40/A gnd NOR3X1_27/C vdd NOR2X1
XNOR2X1_105 INVX1_208/A AND2X2_51/B gnd NOR3X1_21/B vdd NOR2X1
XINVX1_292 dz[12] gnd INVX1_292/Y vdd INVX1
XINVX1_29 vertices[3] gnd INVX1_29/Y vdd INVX1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XINVX1_270 INVX1_270/A gnd INVX1_270/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XNAND2X1_92 AOI22X1_9/A AOI22X1_9/B gnd OAI21X1_97/A vdd NAND2X1
XNAND2X1_70 OAI21X1_52/Y NAND2X1_70/B gnd NAND2X1_70/Y vdd NAND2X1
XNAND2X1_81 OR2X2_9/B OR2X2_9/A gnd NAND3X1_34/B vdd NAND2X1
XAOI21X1_241 INVX1_339/A NAND3X1_456/B NOR2X1_171/Y gnd INVX1_383/A vdd AOI21X1
XFILL_24_1_2 gnd vdd FILL
XAOI21X1_230 NAND3X1_483/B NAND3X1_483/C INVX1_348/Y gnd OAI21X1_461/B vdd AOI21X1
XAOI21X1_252 NAND3X1_528/B INVX1_377/A AND2X2_108/Y gnd NOR3X1_46/B vdd AOI21X1
XAOI21X1_263 OAI21X1_514/Y NAND3X1_543/B OAI21X1_511/Y gnd NOR3X1_52/B vdd AOI21X1
XFILL_7_2_2 gnd vdd FILL
XFILL_15_1_2 gnd vdd FILL
XNAND3X1_201 AOI21X1_83/Y NAND3X1_201/B NAND3X1_201/C gnd NAND3X1_201/Y vdd NAND3X1
XNAND3X1_212 AND2X2_53/B AND2X2_46/Y AOI22X1_25/D gnd AND2X2_53/A vdd NAND3X1
XNAND3X1_223 cos_gamma[5] NAND2X1_70/Y INVX1_198/Y gnd OAI21X1_262/C vdd NAND3X1
XNAND3X1_289 OAI21X1_284/Y OAI21X1_337/C XNOR2X1_34/Y gnd NAND3X1_294/A vdd NAND3X1
XNAND3X1_234 INVX1_207/A OAI21X1_226/Y NAND3X1_234/C gnd NAND3X1_234/Y vdd NAND3X1
XNAND3X1_278 NOR3X1_22/Y INVX1_256/A OAI21X1_251/Y gnd INVX1_224/A vdd NAND3X1
XNAND3X1_267 NAND3X1_267/A NAND3X1_267/B OAI21X1_247/Y gnd NAND3X1_272/A vdd NAND3X1
XNAND3X1_245 INVX1_202/A NAND3X1_248/B OAI21X1_240/Y gnd NAND3X1_251/C vdd NAND3X1
XNAND3X1_256 BUFX2_8/Y OAI21X1_243/C NAND3X1_256/C gnd NAND3X1_259/B vdd NAND3X1
XOAI21X1_408 NOR3X1_42/B NOR3X1_42/C NOR3X1_42/A gnd OAI21X1_408/Y vdd OAI21X1
XFILL_21_1 gnd vdd FILL
XOAI21X1_419 INVX1_259/Y INVX1_18/Y INVX1_299/Y gnd OAI21X1_420/C vdd OAI21X1
XNAND2X1_458 vertices[3] cos_alpha[11] gnd OR2X2_49/B vdd NAND2X1
XNAND2X1_403 AND2X2_91/A AND2X2_91/B gnd NOR3X1_38/A vdd NAND2X1
XNAND2X1_414 NOR2X1_173/A NOR2X1_173/B gnd AOI22X1_45/D vdd NAND2X1
XNAND2X1_425 cos_gamma[14] INVX1_9/A gnd OR2X2_42/B vdd NAND2X1
XNAND2X1_447 NOR2X1_157/Y OAI21X1_500/C gnd INVX1_345/A vdd NAND2X1
XNAND2X1_469 BUFX2_3/Y vertices[14] gnd OAI21X1_450/C vdd NAND2X1
XNAND2X1_436 cos_gamma[10] NAND2X1_70/Y gnd XNOR2X1_80/A vdd NAND2X1
XOAI21X1_68 NOR2X1_47/Y INVX1_72/Y OAI21X1_68/C gnd NOR2X1_57/B vdd OAI21X1
XOAI21X1_57 INVX1_83/A INVX1_84/Y INVX1_69/A gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_13 XNOR2X1_3/B INVX1_25/Y OAI21X1_13/C gnd INVX1_26/A vdd OAI21X1
XOAI21X1_46 INVX1_51/A AND2X2_18/Y NAND3X1_4/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_24 INVX1_1/Y INVX1_50/Y AND2X2_18/A gnd NAND3X1_4/B vdd OAI21X1
XOAI21X1_35 INVX1_36/Y NOR2X1_7/B OAI21X1_64/A gnd OAI21X1_36/C vdd OAI21X1
XOAI21X1_79 OAI21X1_79/A INVX1_105/Y OAI21X1_79/C gnd OAI21X1_79/Y vdd OAI21X1
XOAI21X1_238 OAI21X1_238/A OAI21X1_238/B OAI21X1_238/C gnd OAI21X1_238/Y vdd OAI21X1
XOAI21X1_205 NOR3X1_22/A NOR3X1_22/C NOR3X1_22/B gnd OAI21X1_205/Y vdd OAI21X1
XOAI21X1_249 AOI22X1_29/Y OAI21X1_250/B AND2X2_56/Y gnd OAI21X1_249/Y vdd OAI21X1
XOAI21X1_227 OAI21X1_227/A XNOR2X1_27/Y INVX1_212/A gnd OAI21X1_236/C vdd OAI21X1
XOAI21X1_216 OR2X2_19/A OR2X2_31/B OAI21X1_216/C gnd INVX1_198/A vdd OAI21X1
XAND2X2_49 INVX1_204/Y AND2X2_49/B gnd OR2X2_26/B vdd AND2X2
XNAND2X1_200 OAI21X1_258/C OAI21X1_212/Y gnd OR2X2_23/B vdd NAND2X1
XAND2X2_27 AND2X2_27/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XAND2X2_16 vertices[2] cos_alpha[3] gnd NOR2X1_47/B vdd AND2X2
XAND2X2_38 BUFX2_2/Y vertices[8] gnd NOR2X1_97/B vdd AND2X2
XNAND2X1_211 cos_gamma[1] NAND3X1_399/B gnd OAI21X1_243/C vdd NAND2X1
XNAND2X1_288 INVX1_243/A XOR2X1_19/Y gnd NAND3X1_293/C vdd NAND2X1
XNAND2X1_299 NOR2X1_137/A NOR2X1_137/B gnd NAND3X1_314/C vdd NAND2X1
XNAND2X1_222 OR2X2_26/B OR2X2_26/A gnd INVX1_240/A vdd NAND2X1
XNAND2X1_277 cos_gamma[1] NAND3X1_256/C gnd NOR2X1_137/A vdd NAND2X1
XNAND2X1_233 BUFX2_15/Y vertices[9] gnd INVX1_208/A vdd NAND2X1
XFILL_4_0_2 gnd vdd FILL
XNAND2X1_255 INVX1_254/A NAND3X1_272/B gnd OAI21X1_305/C vdd NAND2X1
XNAND2X1_244 AOI22X1_31/A AOI22X1_31/B gnd NAND3X1_260/C vdd NAND2X1
XNAND2X1_266 INVX1_253/A NAND3X1_268/C gnd OAI21X1_302/C vdd NAND2X1
XFILL_22_2_0 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XNAND3X1_27 OAI21X1_54/Y XOR2X1_6/Y NAND3X1_27/C gnd AND2X2_26/A vdd NAND3X1
XNAND3X1_49 NAND3X1_49/A AOI22X1_9/C AOI22X1_9/D gnd NAND3X1_50/B vdd NAND3X1
XNAND3X1_38 NOR3X1_2/Y NAND3X1_38/B NAND3X1_38/C gnd NAND3X1_59/A vdd NAND3X1
XNAND3X1_16 INVX1_74/A OAI21X1_44/Y OAI21X1_45/Y gnd NAND3X1_19/B vdd NAND3X1
XFILL_27_1_0 gnd vdd FILL
XNAND3X1_405 INVX1_314/A NAND3X1_405/B OAI21X1_387/Y gnd NAND3X1_405/Y vdd NAND3X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_27 dy[3] dx[3] gnd NOR2X1_28/A vdd NOR2X1
XNOR2X1_38 NOR2X1_38/A INVX1_56/Y gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_49 INVX1_68/A NOR2X1_49/B gnd INVX1_79/A vdd NOR2X1
XNOR2X1_16 INVX1_2/Y INVX1_15/Y gnd NOR2X1_16/Y vdd NOR2X1
XNAND3X1_449 NAND3X1_451/B AND2X2_103/A AND2X2_94/Y gnd NAND3X1_450/B vdd NAND3X1
XNAND3X1_438 AOI22X1_55/B OAI21X1_408/Y INVX1_327/Y gnd AOI22X1_47/C vdd NAND3X1
XNAND3X1_416 OAI21X1_389/Y NAND3X1_416/B OAI21X1_399/Y gnd OAI21X1_431/C vdd NAND3X1
XNAND3X1_427 INVX1_359/A INVX1_323/A NAND3X1_429/C gnd NAND3X1_427/Y vdd NAND3X1
XFILL_10_0_0 gnd vdd FILL
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_106 INVX1_211/A NOR2X1_106/B gnd NOR2X1_106/Y vdd NOR2X1
XNOR2X1_139 INVX1_2/Y INVX1_277/Y gnd INVX1_309/A vdd NOR2X1
XNOR2X1_128 NOR2X1_128/A INVX1_251/Y gnd XNOR2X1_36/A vdd NOR2X1
XNOR2X1_117 INVX1_65/Y INVX1_124/Y gnd INVX1_235/A vdd NOR2X1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XINVX1_19 dz[2] gnd INVX1_19/Y vdd INVX1
XINVX1_282 NOR3X1_33/A gnd INVX1_282/Y vdd INVX1
XINVX1_271 INVX1_271/A gnd INVX1_271/Y vdd INVX1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XNAND2X1_71 INVX1_78/Y NOR2X1_48/Y gnd NAND3X1_35/C vdd NAND2X1
XNAND2X1_60 NOR2X1_47/A INVX1_30/A gnd INVX1_77/A vdd NAND2X1
XNAND2X1_93 NAND3X1_47/Y NAND3X1_48/Y gnd NAND3X1_49/A vdd NAND2X1
XNAND2X1_82 XOR2X1_6/B XOR2X1_6/A gnd AND2X2_26/B vdd NAND2X1
XAOI21X1_242 NAND3X1_473/C NAND3X1_473/B INVX1_355/A gnd OAI21X1_482/B vdd AOI21X1
XAOI21X1_264 XNOR2X1_46/Y NAND3X1_494/B OAI21X1_469/B gnd NAND3X1_544/A vdd AOI21X1
XAOI21X1_231 AOI22X1_55/D AOI22X1_55/C NAND3X1_506/B gnd OAI21X1_464/B vdd AOI21X1
XAOI21X1_253 NAND3X1_481/B OAI21X1_458/C NAND3X1_481/C gnd NOR3X1_45/B vdd AOI21X1
XAOI21X1_220 INVX1_308/A AOI22X1_45/D NOR2X1_173/Y gnd OAI21X1_478/A vdd AOI21X1
XNAND3X1_235 NAND3X1_235/A OAI21X1_235/C OAI21X1_232/Y gnd NAND3X1_236/A vdd NAND3X1
XNAND3X1_213 NAND3X1_215/B INVX1_189/Y AND2X2_53/A gnd NAND3X1_214/A vdd NAND3X1
XNAND3X1_202 OAI21X1_219/A NOR2X1_107/A NAND3X1_202/C gnd AOI21X1_98/B vdd NAND3X1
XNAND3X1_246 INVX1_201/Y NAND3X1_251/B NAND3X1_251/C gnd AOI22X1_41/A vdd NAND3X1
XNAND3X1_224 INVX1_200/A AND2X2_61/B NAND3X1_224/C gnd AND2X2_61/A vdd NAND3X1
XNAND3X1_257 BUFX2_9/Y AOI22X1_41/D NAND3X1_257/C gnd NAND3X1_258/C vdd NAND3X1
XNAND3X1_279 cos_gamma[11] INVX1_9/A INVX1_228/Y gnd AND2X2_60/A vdd NAND3X1
XNAND3X1_268 OAI21X1_247/C NAND3X1_268/B NAND3X1_268/C gnd INVX1_254/A vdd NAND3X1
XOAI21X1_409 OAI21X1_410/A NOR3X1_42/Y INVX1_327/Y gnd AOI22X1_46/D vdd OAI21X1
XFILL_21_2 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XNAND2X1_415 dy[13] dx[13] gnd INVX1_325/A vdd NAND2X1
XNAND2X1_426 cos_gamma[13] INVX1_18/A gnd XOR2X1_40/A vdd NAND2X1
XNAND2X1_459 OAI21X1_439/Y OR2X2_49/Y gnd XOR2X1_34/B vdd NAND2X1
XNAND2X1_404 cos_alpha[5] vertices[8] gnd XOR2X1_30/B vdd NAND2X1
XNAND2X1_448 AND2X2_100/B AND2X2_100/A gnd OAI21X1_428/C vdd NAND2X1
XNAND2X1_437 cos_gamma[11] INVX1_43/A gnd OR2X2_44/B vdd NAND2X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_47 OAI21X1_75/B NOR3X1_1/Y OAI21X1_75/A gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_58 INVX1_86/A INVX1_85/Y INVX1_38/Y gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_69 INVX1_16/Y INVX1_46/Y AND2X2_23/Y gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_25 INVX1_52/A OAI21X1_43/C NAND3X1_4/B gnd OAI21X1_26/C vdd OAI21X1
XOAI21X1_14 INVX1_1/Y INVX1_29/Y OAI21X1_7/B gnd AOI21X1_3/A vdd OAI21X1
XOAI21X1_36 OAI21X1_36/A OR2X2_13/B OAI21X1_36/C gnd INVX1_66/A vdd OAI21X1
XOAI21X1_228 INVX1_46/Y INVX1_177/Y NOR2X1_146/A gnd OAI21X1_229/C vdd OAI21X1
XOAI21X1_206 OAI21X1_308/B XOR2X1_12/B OAI21X1_308/C gnd XOR2X1_16/B vdd OAI21X1
XOAI21X1_239 OAI21X1_240/A OAI21X1_240/B INVX1_215/Y gnd OAI21X1_239/Y vdd OAI21X1
XOAI21X1_217 INVX1_65/Y OAI22X1_8/D INVX1_198/A gnd OAI21X1_217/Y vdd OAI21X1
XNAND2X1_223 INVX1_240/A OR2X2_26/Y gnd INVX1_214/A vdd NAND2X1
XNAND2X1_234 INVX1_15/A vertices[8] gnd NOR3X1_21/A vdd NAND2X1
XNAND2X1_201 OR2X2_23/B OR2X2_23/A gnd NAND2X1_202/A vdd NAND2X1
XAND2X2_39 AND2X2_39/A AND2X2_39/B gnd AND2X2_39/Y vdd AND2X2
XAND2X2_28 vertices[3] cos_alpha[4] gnd NOR2X1_77/A vdd AND2X2
XAND2X2_17 INVX1_1/A vertices[5] gnd AND2X2_17/Y vdd AND2X2
XNAND2X1_212 INVX1_199/Y OAI21X1_218/Y gnd AND2X2_61/B vdd NAND2X1
XNAND2X1_289 NAND3X1_285/Y NAND3X1_286/Y gnd NAND3X1_295/C vdd NAND2X1
XNAND2X1_256 cos_gamma[10] INVX1_18/A gnd OAI21X1_314/C vdd NAND2X1
XNAND2X1_267 cos_gamma[3] NAND3X1_457/B gnd OR2X2_31/A vdd NAND2X1
XNAND2X1_245 AOI22X1_41/D NAND3X1_257/C gnd NOR2X1_197/B vdd NAND2X1
XNAND2X1_278 OAI21X1_219/A OAI21X1_219/C gnd NAND2X1_279/B vdd NAND2X1
XFILL_22_2_1 gnd vdd FILL
XOR2X2_50 OR2X2_50/A OR2X2_50/B gnd OR2X2_50/Y vdd OR2X2
XXNOR2X1_1 AND2X2_2/Y XNOR2X1_1/B gnd XNOR2X1_1/Y vdd XNOR2X1
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XAND2X2_1 OR2X2_1/Y AND2X2_1/B gnd NOR2X1_5/B vdd AND2X2
XNOR2X1_28 NOR2X1_28/A INVX1_33/Y gnd XNOR2X1_7/A vdd NOR2X1
XNAND3X1_28 OAI21X1_39/Y AND2X2_26/A NAND3X1_28/C gnd INVX1_84/A vdd NAND3X1
XNAND3X1_39 INVX1_99/Y OAI22X1_4/Y NAND3X1_47/C gnd AOI22X1_9/A vdd NAND3X1
XNOR2X1_17 NOR2X1_17/A AND2X2_5/Y gnd NOR2X1_18/A vdd NOR2X1
XNAND3X1_17 INVX1_74/Y AOI22X1_7/D AOI22X1_3/D gnd NAND3X1_19/A vdd NAND3X1
XNAND3X1_406 OAI21X1_432/C NAND3X1_406/B INVX1_313/Y gnd NAND3X1_407/B vdd NAND3X1
XFILL_27_1_1 gnd vdd FILL
XNAND3X1_417 OAI21X1_431/C OAI21X1_401/Y INVX1_315/Y gnd NAND3X1_418/B vdd NAND3X1
XNAND3X1_439 AOI22X1_47/C AOI22X1_47/D NAND3X1_439/C gnd NAND3X1_443/B vdd NAND3X1
XNAND3X1_428 BUFX2_5/Y NOR2X1_173/A NAND3X1_432/C gnd NAND3X1_431/B vdd NAND3X1
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_39 INVX1_40/Y NOR2X1_39/B gnd NOR2X1_40/A vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_118 INVX1_2/Y INVX1_241/Y gnd XOR2X1_17/B vdd NOR2X1
XFILL_18_1_1 gnd vdd FILL
XNOR2X1_129 XNOR2X1_23/A XOR2X1_12/A gnd NOR2X1_129/Y vdd NOR2X1
XNOR2X1_107 NOR2X1_107/A NOR2X1_107/B gnd NOR2X1_107/Y vdd NOR2X1
XINVX1_250 dz[11] gnd INVX1_250/Y vdd INVX1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XINVX1_294 XOR2X1_24/Y gnd INVX1_294/Y vdd INVX1
XINVX1_283 INVX1_283/A gnd OR2X2_33/B vdd INVX1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XNAND2X1_50 NAND2X1_50/A OR2X2_7/Y gnd NOR2X1_39/B vdd NAND2X1
XNAND2X1_61 NOR2X1_47/A NOR2X1_47/B gnd OAI21X1_68/C vdd NAND2X1
XNAND2X1_94 OAI21X1_53/Y NAND3X1_35/C gnd OAI22X1_8/D vdd NAND2X1
XNAND2X1_83 INVX1_78/A NOR2X1_48/B gnd NAND3X1_57/C vdd NAND2X1
XNAND2X1_72 dy[5] dx[5] gnd INVX1_81/A vdd NAND2X1
XAOI21X1_265 NAND3X1_545/C NAND3X1_545/B INVX1_384/Y gnd OAI21X1_518/A vdd AOI21X1
XAOI21X1_221 NAND3X1_470/A NAND3X1_470/B OAI21X1_497/B gnd NOR3X1_44/C vdd AOI21X1
XAOI21X1_243 XOR2X1_34/A INVX1_371/Y NOR2X1_181/Y gnd XOR2X1_44/B vdd AOI21X1
XAOI21X1_232 AOI22X1_54/D AOI22X1_54/C NAND3X1_506/B gnd OAI21X1_479/A vdd AOI21X1
XAOI21X1_210 OAI21X1_348/Y INVX1_276/Y NOR3X1_35/Y gnd NAND3X1_424/A vdd AOI21X1
XAOI21X1_254 OAI21X1_499/Y OAI21X1_500/Y NOR2X1_196/Y gnd OAI21X1_504/A vdd AOI21X1
XNAND3X1_236 NAND3X1_236/A OAI21X1_236/Y OAI21X1_271/B gnd NAND3X1_240/C vdd NAND3X1
XNAND3X1_203 OAI21X1_219/A NOR2X1_107/A NOR2X1_107/B gnd NAND3X1_204/B vdd NAND3X1
XNAND3X1_214 NAND3X1_214/A NAND3X1_214/B OAI21X1_201/Y gnd NAND3X1_217/B vdd NAND3X1
XNAND3X1_269 INVX1_254/A AOI22X1_29/D AND2X2_55/Y gnd NAND3X1_272/B vdd NAND3X1
XNAND3X1_225 INVX1_200/Y NAND3X1_225/B NAND3X1_225/C gnd AND2X2_54/B vdd NAND3X1
XNAND3X1_247 INVX1_202/A INVX1_248/A OAI21X1_239/Y gnd NAND3X1_252/B vdd NAND3X1
XNAND3X1_258 cos_gamma[1] NAND3X1_399/B NAND3X1_258/C gnd NAND3X1_259/C vdd NAND3X1
XNAND2X1_416 AOI22X1_46/A AOI22X1_46/B gnd NAND3X1_439/C vdd NAND2X1
XNAND2X1_405 cos_alpha[4] vertices[9] gnd XOR2X1_29/A vdd NAND2X1
XNAND2X1_427 OR2X2_42/B OR2X2_42/A gnd NAND2X1_428/A vdd NAND2X1
XNAND2X1_449 OAI21X1_478/A AND2X2_100/Y gnd NAND3X1_459/B vdd NAND2X1
XNAND2X1_438 cos_gamma[6] NAND3X1_457/B gnd NAND2X1_439/B vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_48 NOR2X1_46/Y NOR2X1_47/Y INVX1_72/A gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_59 INVX1_38/Y INVX1_86/A INVX1_85/A gnd INVX1_90/A vdd OAI21X1
XOAI21X1_26 INVX1_16/Y INVX1_15/Y OAI21X1_26/C gnd NAND3X1_5/B vdd OAI21X1
XOAI21X1_15 OR2X2_3/B AND2X2_18/A AOI21X1_3/A gnd XNOR2X1_4/A vdd OAI21X1
XOAI21X1_37 INVX1_65/Y INVX1_9/Y INVX1_66/A gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_229 OAI21X1_229/A OAI21X1_277/C OAI21X1_229/C gnd XOR2X1_14/A vdd OAI21X1
XAND2X2_18 AND2X2_18/A INVX1_102/A gnd AND2X2_18/Y vdd AND2X2
XOAI21X1_207 INVX1_139/Y OAI21X1_207/B AND2X2_57/B gnd AOI22X1_38/A vdd OAI21X1
XAND2X2_29 cos_alpha[3] vertices[4] gnd NOR2X1_77/B vdd AND2X2
XOAI21X1_218 OAI21X1_218/A OAI21X1_243/C AND2X2_48/A gnd OAI21X1_218/Y vdd OAI21X1
XNAND2X1_224 vertices[2] cos_alpha[8] gnd XOR2X1_13/B vdd NAND2X1
XNAND2X1_235 BUFX2_2/Y vertices[10] gnd AND2X2_51/B vdd NAND2X1
XNAND2X1_257 cos_gamma[7] NAND2X1_70/Y gnd NOR2X1_133/A vdd NAND2X1
XNAND2X1_268 OR2X2_31/B OR2X2_31/A gnd OAI21X1_263/C vdd NAND2X1
XNAND2X1_202 NAND2X1_202/A OR2X2_23/Y gnd OR2X2_24/A vdd NAND2X1
XNAND2X1_246 dy[10] dx[10] gnd INVX1_219/A vdd NAND2X1
XNAND2X1_213 INVX1_199/A AND2X2_48/Y gnd NAND3X1_224/C vdd NAND2X1
XNAND2X1_279 NAND3X1_199/Y NAND2X1_279/B gnd AOI22X1_32/C vdd NAND2X1
XFILL_22_2_2 gnd vdd FILL
XOR2X2_51 OR2X2_51/A OR2X2_51/B gnd OR2X2_51/Y vdd OR2X2
XOR2X2_40 OR2X2_40/A OR2X2_40/B gnd OR2X2_40/Y vdd OR2X2
XXNOR2X1_2 XNOR2X1_2/A INVX1_19/Y gnd OR2X2_4/B vdd XNOR2X1
XFILL_13_2_2 gnd vdd FILL
XINVX1_2 vertices[0] gnd INVX1_2/Y vdd INVX1
XOAI21X1_390 OR2X2_33/B OR2X2_33/A OR2X2_32/Y gnd INVX1_317/A vdd OAI21X1
XAND2X2_2 OR2X2_2/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XFILL_27_1_2 gnd vdd FILL
XNAND3X1_29 INVX1_69/Y INVX1_84/A INVX1_83/Y gnd NAND3X1_30/C vdd NAND3X1
XNAND3X1_18 OAI21X1_68/C OAI21X1_41/Y INVX1_72/Y gnd NAND3X1_18/Y vdd NAND3X1
XNOR2X1_29 INVX1_21/A XNOR2X1_9/Y gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_18 NOR2X1_18/A INVX1_17/Y gnd INVX1_18/A vdd NOR2X1
XNAND3X1_407 INVX1_314/Y NAND3X1_407/B OAI21X1_388/Y gnd NAND3X1_407/Y vdd NAND3X1
XNAND3X1_418 OAI21X1_380/Y NAND3X1_418/B OAI21X1_402/Y gnd OAI21X1_430/C vdd NAND3X1
XNAND3X1_429 INVX1_359/A INVX1_323/Y NAND3X1_429/C gnd NAND3X1_508/B vdd NAND3X1
XFILL_2_1_2 gnd vdd FILL
XFILL_10_0_2 gnd vdd FILL
XNOR2X1_119 INVX1_204/Y XOR2X1_17/Y gnd INVX1_242/A vdd NOR2X1
XFILL_18_1_2 gnd vdd FILL
XNOR2X1_108 dy[10] dx[10] gnd NOR2X1_109/A vdd NOR2X1
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XINVX1_262 INVX1_262/A gnd INVX1_262/Y vdd INVX1
XINVX1_284 NOR3X1_26/A gnd INVX1_284/Y vdd INVX1
XINVX1_273 INVX1_273/A gnd INVX1_273/Y vdd INVX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XNAND2X1_73 OAI21X1_54/Y NAND3X1_27/C gnd OAI21X1_66/B vdd NAND2X1
XNAND2X1_95 dy[6] dx[6] gnd INVX1_107/A vdd NAND2X1
XNAND2X1_51 INVX1_40/Y NOR2X1_39/B gnd INVX1_58/A vdd NAND2X1
XNAND2X1_62 vertices[2] cos_alpha[3] gnd NOR2X1_46/B vdd NAND2X1
XNAND2X1_40 vertices[2] BUFX2_12/Y gnd INVX1_51/A vdd NAND2X1
XNAND2X1_84 vertices[0] cos_alpha[6] gnd INVX1_97/A vdd NAND2X1
XAOI21X1_200 AND2X2_77/Y OAI21X1_343/Y NOR3X1_29/C gnd NOR3X1_37/A vdd AOI21X1
XAOI22X1_60 AOI22X1_60/A AOI22X1_60/B AOI22X1_60/C AOI22X1_60/D gnd NOR3X1_52/C vdd
+ AOI22X1
XAOI21X1_266 INVX1_330/Y OAI21X1_470/Y INVX1_385/Y gnd OAI21X1_518/C vdd AOI21X1
XAOI21X1_244 AOI22X1_58/A AOI22X1_58/B INVX1_373/A gnd OAI22X1_12/C vdd AOI21X1
XAOI21X1_255 NAND3X1_533/A NAND3X1_533/B NAND3X1_533/C gnd NOR3X1_47/C vdd AOI21X1
XAOI21X1_222 NAND3X1_472/Y NAND3X1_474/Y INVX1_357/A gnd OAI21X1_456/A vdd AOI21X1
XAOI21X1_233 OAI21X1_465/Y OAI21X1_464/Y INVX1_341/A gnd OAI21X1_467/A vdd AOI21X1
XAOI21X1_211 NAND2X1_351/B NAND2X1_351/A INVX1_8/Y gnd NAND3X1_432/B vdd AOI21X1
XNAND3X1_226 INVX1_207/A NAND3X1_233/A OAI21X1_225/Y gnd NAND3X1_226/Y vdd NAND3X1
XNAND3X1_237 INVX1_246/A OAI21X1_235/Y NAND3X1_237/C gnd NAND3X1_240/B vdd NAND3X1
XNAND3X1_204 INVX1_7/A NAND3X1_204/B NAND3X1_204/C gnd NAND3X1_204/Y vdd NAND3X1
XNAND3X1_215 INVX1_189/A NAND3X1_215/B AND2X2_53/A gnd AND2X2_56/B vdd NAND3X1
XNAND3X1_248 INVX1_202/Y NAND3X1_248/B OAI21X1_240/Y gnd NAND3X1_252/C vdd NAND3X1
XNAND3X1_259 INVX1_217/A NAND3X1_259/B NAND3X1_259/C gnd NAND3X1_261/B vdd NAND3X1
XNAND2X1_417 AOI22X1_47/A AOI22X1_47/B gnd NAND3X1_440/C vdd NAND2X1
XNAND2X1_428 NAND2X1_428/A OR2X2_42/Y gnd OR2X2_43/B vdd NAND2X1
XNAND2X1_406 cos_alpha[3] vertices[10] gnd OR2X2_57/A vdd NAND2X1
XNAND2X1_439 NOR2X1_166/B NAND2X1_439/B gnd INVX1_337/A vdd NAND2X1
XFILL_7_0_2 gnd vdd FILL
XOAI21X1_16 INVX1_2/Y INVX1_28/Y AND2X2_9/A gnd NAND3X1_3/C vdd OAI21X1
XOAI21X1_27 NOR3X1_2/A NOR3X1_2/C INVX1_44/Y gnd NAND3X1_8/A vdd OAI21X1
XOAI21X1_49 NOR3X1_1/B NOR3X1_1/C NOR3X1_1/A gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_38 NOR2X1_43/A INVX1_37/Y OAI21X1_38/C gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_208 OR2X2_17/B OR2X2_17/A AOI22X1_30/A gnd INVX1_223/A vdd OAI21X1
XOAI21X1_219 OAI21X1_219/A OAI21X1_219/B OAI21X1_219/C gnd OAI21X1_242/A vdd OAI21X1
XAND2X2_19 AND2X2_19/A OR2X2_8/Y gnd NOR2X1_53/B vdd AND2X2
XNAND2X1_225 vertices[4] cos_alpha[7] gnd OAI21X1_272/C vdd NAND2X1
XNAND2X1_258 INVX1_230/A NOR2X1_115/Y gnd OAI21X1_316/C vdd NAND2X1
XNAND2X1_236 AND2X2_44/Y AND2X2_52/Y gnd OAI21X1_279/C vdd NAND2X1
XNAND2X1_269 cos_gamma[4] NAND3X1_457/B gnd OR2X2_37/B vdd NAND2X1
XNAND2X1_203 OR2X2_24/B OR2X2_24/A gnd AND2X2_58/B vdd NAND2X1
XNAND2X1_214 INVX1_199/Y AND2X2_48/Y gnd NAND3X1_225/C vdd NAND2X1
XNAND2X1_247 NAND3X1_261/B NAND3X1_261/C gnd OAI21X1_265/B vdd NAND2X1
XFILL_25_2_0 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XOR2X2_41 OR2X2_41/A OR2X2_41/B gnd OR2X2_41/Y vdd OR2X2
XOR2X2_52 OR2X2_52/A OR2X2_52/B gnd OR2X2_52/Y vdd OR2X2
XOR2X2_30 OR2X2_30/A OR2X2_30/B gnd OR2X2_30/Y vdd OR2X2
XOR2X2_1 OR2X2_1/A dz[0] gnd OR2X2_1/Y vdd OR2X2
XXNOR2X1_3 XOR2X1_1/Y XNOR2X1_3/B gnd XOR2X1_2/A vdd XNOR2X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_22_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XOAI21X1_380 NOR3X1_33/A NOR3X1_33/B OAI21X1_380/C gnd OAI21X1_380/Y vdd OAI21X1
XOAI21X1_391 INVX1_177/Y INVX1_146/Y OAI21X1_484/A gnd OAI21X1_392/C vdd OAI21X1
XAND2X2_3 INVX1_14/Y AND2X2_3/B gnd AND2X2_4/A vdd AND2X2
XNAND3X1_19 NAND3X1_19/A NAND3X1_19/B OAI21X1_46/Y gnd OAI21X1_75/C vdd NAND3X1
XNOR2X1_19 dy[2] dx[2] gnd NOR2X1_20/A vdd NOR2X1
XNAND3X1_419 INVX1_322/A OAI21X1_430/C OAI21X1_403/Y gnd NAND3X1_424/B vdd NAND3X1
XNAND3X1_408 INVX1_317/A NAND3X1_408/B NAND3X1_408/C gnd AND2X2_91/A vdd NAND3X1
XNOR2X1_109 NOR2X1_109/A INVX1_219/Y gnd XNOR2X1_33/A vdd NOR2X1
XINVX1_241 cos_alpha[11] gnd INVX1_241/Y vdd INVX1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XINVX1_285 INVX1_285/A gnd INVX1_285/Y vdd INVX1
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XINVX1_274 INVX1_274/A gnd INVX1_274/Y vdd INVX1
XINVX1_252 XOR2X1_21/Y gnd NOR3X1_25/A vdd INVX1
XNAND2X1_63 NAND3X1_15/Y OAI21X1_42/Y gnd OAI21X1_75/A vdd NAND2X1
XNAND2X1_96 INVX1_118/A OAI21X1_83/Y gnd NAND2X1_97/B vdd NAND2X1
XNAND2X1_74 INVX1_82/Y OAI21X1_66/B gnd NAND3X1_28/C vdd NAND2X1
XNAND2X1_85 INVX1_97/Y NOR2X1_57/B gnd INVX1_98/A vdd NAND2X1
XNAND2X1_52 INVX1_39/Y NOR2X1_40/Y gnd NAND3X1_9/B vdd NAND2X1
XNAND2X1_41 AOI22X1_2/B INVX1_52/Y gnd NAND3X1_4/C vdd NAND2X1
XNAND2X1_30 OR2X2_6/B OR2X2_6/A gnd AOI21X1_1/B vdd NAND2X1
XAOI21X1_234 OAI21X1_462/Y OAI21X1_463/Y INVX1_341/Y gnd OAI21X1_467/B vdd AOI21X1
XAOI21X1_223 NAND3X1_475/Y NAND3X1_476/Y INVX1_357/Y gnd OAI21X1_456/B vdd AOI21X1
XAOI21X1_201 NAND3X1_413/C INVX1_320/A XNOR2X1_44/Y gnd NOR3X1_37/B vdd AOI21X1
XAOI21X1_212 NAND3X1_431/C NAND3X1_431/B INVX1_308/Y gnd NOR3X1_42/C vdd AOI21X1
XAOI21X1_245 AOI22X1_57/A AOI22X1_57/B INVX1_373/Y gnd OAI22X1_12/D vdd AOI21X1
XAOI21X1_256 NAND3X1_532/A NAND3X1_532/B NAND3X1_532/C gnd NOR3X1_47/B vdd AOI21X1
XAOI22X1_50 OR2X2_35/Y AOI22X1_50/B AOI22X1_50/C AOI22X1_50/D gnd AOI22X1_50/Y vdd
+ AOI22X1
XNAND3X1_205 INVX1_184/A NAND3X1_205/B NAND3X1_205/C gnd NAND3X1_208/C vdd NAND3X1
XNAND3X1_227 OAI21X1_226/Y INVX1_207/Y NAND3X1_234/C gnd NAND3X1_227/Y vdd NAND3X1
XNAND3X1_216 AND2X2_56/B AOI22X1_26/D AND2X2_47/Y gnd AND2X2_56/A vdd NAND3X1
XNAND3X1_249 INVX1_201/A NAND3X1_252/B NAND3X1_252/C gnd NAND3X1_254/C vdd NAND3X1
XNAND3X1_238 NAND3X1_240/B NAND3X1_240/C OAI21X1_238/C gnd NAND3X1_239/B vdd NAND3X1
XOAI22X1_1 INVX1_8/Y INVX1_9/Y INVX1_7/Y NOR2X1_7/B gnd OAI22X1_1/Y vdd OAI22X1
XNAND2X1_418 INVX1_303/A XNOR2X1_42/Y gnd AOI22X1_49/A vdd NAND2X1
XNAND2X1_429 OR2X2_43/B OR2X2_43/A gnd NAND2X1_430/A vdd NAND2X1
XNAND2X1_407 BUFX2_2/Y vertices[13] gnd OR2X2_40/B vdd NAND2X1
XOAI21X1_39 OR2X2_7/B OR2X2_7/A OAI21X1_39/C gnd OAI21X1_39/Y vdd OAI21X1
XOAI21X1_28 INVX1_67/A INVX1_68/A OAI22X1_3/Y gnd XNOR2X1_11/A vdd OAI21X1
XOAI21X1_17 NOR2X1_25/A AND2X2_8/Y INVX1_30/A gnd INVX1_31/A vdd OAI21X1
XOAI21X1_209 OAI22X1_8/A INVX1_9/Y OAI21X1_311/A gnd OAI21X1_210/C vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XNAND2X1_259 INVX1_232/A NOR2X1_116/Y gnd NAND2X1_260/B vdd NAND2X1
XNAND2X1_226 vertices[4] cos_alpha[6] gnd NOR2X1_142/A vdd NAND2X1
XNAND2X1_237 NAND3X1_232/A OAI21X1_230/Y gnd NOR2X1_106/B vdd NAND2X1
XNAND2X1_215 INVX1_199/A OAI21X1_218/Y gnd NAND3X1_225/B vdd NAND2X1
XNAND2X1_204 AND2X2_58/B OR2X2_24/Y gnd XNOR2X1_31/B vdd NAND2X1
XNAND2X1_248 INVX1_220/Y OAI21X1_265/B gnd NAND3X1_263/C vdd NAND2X1
XFILL_25_2_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XOR2X2_53 OR2X2_53/A OR2X2_53/B gnd OR2X2_53/Y vdd OR2X2
XOR2X2_42 OR2X2_42/A OR2X2_42/B gnd OR2X2_42/Y vdd OR2X2
XOR2X2_31 OR2X2_31/A OR2X2_31/B gnd OR2X2_31/Y vdd OR2X2
XOR2X2_2 OR2X2_2/A dz[1] gnd OR2X2_2/Y vdd OR2X2
XXNOR2X1_4 XNOR2X1_4/A INVX1_48/A gnd AND2X2_8/A vdd XNOR2X1
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XINVX1_4 dy[0] gnd INVX1_4/Y vdd INVX1
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_381 INVX1_2/Y INVX1_310/Y OAI21X1_491/A gnd OAI21X1_382/C vdd OAI21X1
XOAI21X1_392 OR2X2_32/B OAI21X1_443/C OAI21X1_392/C gnd OR2X2_39/A vdd OAI21X1
XOAI21X1_370 OAI22X1_8/A INVX1_43/Y OAI21X1_476/A gnd AND2X2_85/B vdd OAI21X1
XAND2X2_4 AND2X2_4/A INVX1_6/Y gnd AND2X2_4/Y vdd AND2X2
XNAND3X1_409 INVX1_317/Y NAND3X1_409/B NAND3X1_409/C gnd AND2X2_91/B vdd NAND3X1
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XINVX1_264 INVX1_264/A gnd INVX1_264/Y vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XINVX1_275 XOR2X1_18/B gnd INVX1_275/Y vdd INVX1
XINVX1_220 XOR2X1_15/Y gnd INVX1_220/Y vdd INVX1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XNAND2X1_97 INVX1_110/Y NAND2X1_97/B gnd NAND3X1_66/C vdd NAND2X1
XNAND2X1_20 NAND2X1_20/A NAND2X1_20/B gnd XNOR2X1_9/B vdd NAND2X1
XNAND2X1_75 NAND3X1_32/B OAI21X1_58/Y gnd NAND2X1_76/B vdd NAND2X1
XNAND2X1_42 NAND3X1_5/A NAND3X1_5/B gnd NAND2X1_43/B vdd NAND2X1
XNAND2X1_31 XNOR2X1_9/B XOR2X1_4/Y gnd INVX1_61/A vdd NAND2X1
XNAND2X1_86 vertices[1] cos_alpha[5] gnd INVX1_99/A vdd NAND2X1
XNAND2X1_64 AOI22X1_2/B AND2X2_17/Y gnd AOI22X1_3/D vdd NAND2X1
XNAND2X1_53 cos_gamma[3] INVX1_18/A gnd OAI21X1_64/A vdd NAND2X1
XAOI21X1_246 OAI22X1_12/Y NAND3X1_518/B INVX1_376/Y gnd OAI21X1_495/A vdd AOI21X1
XAOI21X1_257 NAND3X1_535/B NAND3X1_535/A AND2X2_109/Y gnd NOR3X1_49/B vdd AOI21X1
XAOI21X1_235 NAND3X1_498/C OAI21X1_467/Y AND2X2_102/Y gnd OAI21X1_469/B vdd AOI21X1
XAOI21X1_224 NAND3X1_472/Y NAND3X1_474/Y INVX1_357/Y gnd OR2X2_58/A vdd AOI21X1
XAOI21X1_213 NAND3X1_434/B NAND3X1_434/C XOR2X1_31/Y gnd OAI21X1_410/A vdd AOI21X1
XAOI21X1_202 OAI21X1_396/Y NAND3X1_411/B OAI21X1_395/Y gnd NOR3X1_36/A vdd AOI21X1
XAOI22X1_51 OR2X2_41/Y AOI22X1_51/B AOI22X1_51/C AOI22X1_51/D gnd AOI22X1_51/Y vdd
+ AOI22X1
XAOI22X1_40 INVX1_1/A vertices[12] INVX1_10/A vertices[11] gnd NOR3X1_27/B vdd AOI22X1
XNAND3X1_228 INVX1_209/Y OAI21X1_231/Y OAI21X1_279/C gnd NAND3X1_232/A vdd NAND3X1
XNAND3X1_217 INVX1_190/A NAND3X1_217/B AND2X2_56/A gnd AND2X2_57/B vdd NAND3X1
XNAND3X1_206 BUFX2_7/Y INVX1_171/A NAND3X1_399/B gnd AND2X2_48/B vdd NAND3X1
XNAND3X1_239 INVX1_214/A NAND3X1_239/B OAI21X1_237/Y gnd NAND3X1_244/A vdd NAND3X1
XOAI22X1_2 INVX1_2/Y INVX1_46/Y INVX1_45/Y INVX1_28/Y gnd OAI22X1_2/Y vdd OAI22X1
XNAND2X1_419 INVX1_303/Y OAI21X1_418/B gnd AOI22X1_49/B vdd NAND2X1
XNAND2X1_408 NAND3X1_411/B OAI21X1_396/Y gnd NAND3X1_412/C vdd NAND2X1
XOAI21X1_29 INVX1_32/Y NOR2X1_28/A INVX1_33/A gnd XOR2X1_5/B vdd OAI21X1
XOAI21X1_18 INVX1_31/Y AND2X2_9/Y INVX1_17/Y gnd NAND3X1_8/C vdd OAI21X1
XFILL_12_2 gnd vdd FILL
XNAND2X1_216 XOR2X1_11/B XOR2X1_11/A gnd NAND2X1_217/A vdd NAND2X1
XNAND2X1_205 OR2X2_25/B OR2X2_25/A gnd AND2X2_59/A vdd NAND2X1
XNAND2X1_227 OAI22X1_7/Y XOR2X1_13/Y gnd NAND3X1_233/A vdd NAND2X1
XNAND2X1_238 NAND3X1_234/Y NAND3X1_233/Y gnd OAI21X1_271/B vdd NAND2X1
XNAND2X1_249 AND2X2_61/A AND2X2_54/B gnd NAND3X1_264/B vdd NAND2X1
XFILL_25_2_2 gnd vdd FILL
XFILL_0_2_2 gnd vdd FILL
XFILL_16_2_2 gnd vdd FILL
XOR2X2_32 OR2X2_32/A OR2X2_32/B gnd OR2X2_32/Y vdd OR2X2
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XOR2X2_54 OR2X2_54/A OR2X2_54/B gnd OR2X2_54/Y vdd OR2X2
XOR2X2_43 OR2X2_43/A OR2X2_43/B gnd OR2X2_43/Y vdd OR2X2
XXNOR2X1_5 INVX1_67/A XNOR2X1_5/B gnd XNOR2X1_6/A vdd XNOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 dx[0] gnd INVX1_5/Y vdd INVX1
.ends

