magic
tech scmos
magscale 1 2
timestamp 1651764895
<< metal1 >>
rect 3112 5806 3118 5814
rect 3126 5806 3132 5814
rect 3140 5806 3146 5814
rect 3154 5806 3160 5814
rect 1288 5776 1292 5784
rect 132 5757 147 5763
rect 964 5756 972 5764
rect 1140 5756 1148 5764
rect 1540 5757 1596 5763
rect 109 5737 124 5743
rect 372 5737 387 5743
rect 285 5717 323 5723
rect 525 5717 540 5723
rect 669 5723 675 5736
rect 596 5717 627 5723
rect 637 5717 675 5723
rect 765 5723 771 5743
rect 765 5717 803 5723
rect 1005 5723 1011 5743
rect 1204 5737 1235 5743
rect 1645 5737 1699 5743
rect 1940 5737 1964 5743
rect 2525 5737 2540 5743
rect 2724 5737 2739 5743
rect 3028 5737 3043 5743
rect 3501 5743 3507 5763
rect 3540 5756 3548 5764
rect 4180 5757 4204 5763
rect 4509 5757 4540 5763
rect 4765 5757 4787 5763
rect 3300 5737 3315 5743
rect 973 5717 1011 5723
rect 1060 5717 1091 5723
rect 1357 5717 1388 5723
rect 1453 5717 1491 5723
rect 1629 5717 1644 5723
rect 1917 5717 1932 5723
rect 2557 5717 2572 5723
rect 3389 5723 3395 5743
rect 3501 5737 3516 5743
rect 3677 5737 3715 5743
rect 3812 5737 3827 5743
rect 3901 5737 3955 5743
rect 4045 5737 4083 5743
rect 4132 5737 4163 5743
rect 4333 5737 4387 5743
rect 4573 5743 4579 5756
rect 4452 5737 4467 5743
rect 4557 5737 4579 5743
rect 4749 5737 4764 5743
rect 4781 5743 4787 5757
rect 5517 5757 5548 5763
rect 4781 5737 4803 5743
rect 4941 5737 4972 5743
rect 5341 5737 5395 5743
rect 5581 5743 5587 5756
rect 5460 5737 5475 5743
rect 5565 5737 5587 5743
rect 3341 5717 3379 5723
rect 3389 5717 3412 5723
rect 3341 5704 3347 5717
rect 3404 5712 3412 5717
rect 3485 5717 3516 5723
rect 3533 5717 3571 5723
rect 404 5697 419 5703
rect 1556 5697 1619 5703
rect 2488 5696 2492 5704
rect 2637 5697 2652 5703
rect 2984 5696 2988 5704
rect 3565 5697 3571 5717
rect 3645 5717 3667 5723
rect 3940 5717 3987 5723
rect 4093 5717 4115 5723
rect 4173 5717 4188 5723
rect 4477 5717 4499 5723
rect 4516 5717 4547 5723
rect 4612 5717 4684 5723
rect 4740 5717 4819 5723
rect 5485 5717 5507 5723
rect 5524 5717 5555 5723
rect 5885 5717 5916 5723
rect 6052 5717 6067 5723
rect 4189 5697 4195 5716
rect 5197 5697 5219 5703
rect 429 5677 483 5683
rect 1997 5677 2028 5683
rect 2845 5677 2899 5683
rect 3396 5677 3443 5683
rect 4820 5676 4822 5684
rect 324 5656 326 5664
rect 728 5636 732 5644
rect 1028 5636 1030 5644
rect 1450 5636 1452 5644
rect 2164 5636 2166 5644
rect 2228 5636 2230 5644
rect 3748 5636 3752 5644
rect 3882 5636 3884 5644
rect 4404 5636 4406 5644
rect 5172 5636 5174 5644
rect 5284 5636 5288 5644
rect 5412 5636 5414 5644
rect 6218 5636 6220 5644
rect 1560 5606 1566 5614
rect 1574 5606 1580 5614
rect 1588 5606 1594 5614
rect 1602 5606 1608 5614
rect 4632 5606 4638 5614
rect 4646 5606 4652 5614
rect 4660 5606 4666 5614
rect 4674 5606 4680 5614
rect 148 5576 150 5584
rect 1300 5576 1302 5584
rect 4554 5576 4556 5584
rect 4804 5576 4808 5584
rect 5594 5556 5596 5564
rect 5940 5556 5942 5564
rect 234 5536 236 5544
rect 4612 5536 4614 5544
rect 5300 5536 5302 5544
rect 5676 5537 5731 5543
rect 1757 5504 1763 5523
rect 2237 5517 2259 5523
rect 2292 5517 2307 5523
rect 2797 5517 2851 5523
rect 3917 5517 3932 5523
rect 4461 5517 4492 5523
rect 5325 5517 5340 5523
rect 29 5497 44 5503
rect 829 5497 851 5503
rect 996 5497 1027 5503
rect 1108 5497 1123 5503
rect 1764 5497 1827 5503
rect 1924 5497 1955 5503
rect 1965 5497 2019 5503
rect 2733 5497 2748 5503
rect 3053 5497 3091 5503
rect 4029 5497 4044 5503
rect 4340 5497 4419 5503
rect 4509 5497 4547 5503
rect 5220 5497 5299 5503
rect 5604 5497 5651 5503
rect 5853 5503 5859 5523
rect 6029 5517 6051 5523
rect 5821 5497 5859 5503
rect 5885 5497 5916 5503
rect 5949 5497 5987 5503
rect 6221 5497 6236 5503
rect 452 5477 483 5483
rect 909 5483 915 5496
rect 804 5477 819 5483
rect 893 5477 915 5483
rect 1053 5477 1075 5483
rect 1149 5477 1171 5483
rect 1149 5464 1155 5477
rect 2077 5477 2092 5483
rect 2660 5477 2684 5483
rect 2740 5477 2755 5483
rect 3117 5477 3180 5483
rect 3260 5477 3276 5483
rect 3260 5476 3268 5477
rect 3581 5477 3596 5483
rect 3949 5477 3980 5483
rect 4164 5477 4179 5483
rect 4349 5477 4364 5483
rect 4372 5477 4403 5483
rect 5236 5477 5283 5483
rect 5620 5477 5635 5483
rect 5736 5477 5763 5483
rect 5773 5477 5788 5483
rect 6205 5477 6252 5483
rect 916 5457 931 5463
rect 948 5457 979 5463
rect 1092 5457 1116 5463
rect 1549 5457 1635 5463
rect 2013 5457 2035 5463
rect 2708 5456 2716 5464
rect 4148 5456 4156 5464
rect 5956 5457 5971 5463
rect 548 5436 552 5444
rect 1466 5436 1468 5444
rect 1684 5436 1686 5444
rect 2266 5436 2268 5444
rect 2314 5436 2316 5444
rect 2504 5436 2508 5444
rect 3332 5436 3334 5444
rect 3629 5437 3644 5443
rect 3812 5436 3816 5444
rect 3112 5406 3118 5414
rect 3126 5406 3132 5414
rect 3140 5406 3146 5414
rect 3154 5406 3160 5414
rect 660 5376 664 5384
rect 772 5376 776 5384
rect 1000 5376 1004 5384
rect 2077 5377 2092 5383
rect 2296 5376 2300 5384
rect 2424 5376 2428 5384
rect 3592 5376 3596 5384
rect 3933 5377 3948 5383
rect 4018 5377 4060 5383
rect 4093 5377 4108 5383
rect 5124 5377 5139 5383
rect 5914 5376 5916 5384
rect 6202 5376 6204 5384
rect 237 5357 259 5363
rect 500 5356 508 5364
rect 925 5344 931 5363
rect 3956 5357 3971 5363
rect 68 5337 115 5343
rect 285 5337 332 5343
rect 365 5337 419 5343
rect 532 5337 547 5343
rect 541 5324 547 5337
rect 717 5337 732 5343
rect 852 5337 867 5343
rect 877 5337 915 5343
rect 932 5337 947 5343
rect 1524 5337 1555 5343
rect 1700 5337 1715 5343
rect 2040 5336 2044 5344
rect 2461 5337 2508 5343
rect 2573 5337 2620 5343
rect 3085 5337 3171 5343
rect 3348 5337 3379 5343
rect 3524 5337 3539 5343
rect 77 5317 92 5323
rect 301 5317 316 5323
rect 381 5317 396 5323
rect 1076 5317 1107 5323
rect 1197 5323 1203 5336
rect 3629 5324 3635 5343
rect 4173 5337 4204 5343
rect 4253 5337 4284 5343
rect 4445 5343 4451 5363
rect 5373 5357 5395 5363
rect 5844 5356 5852 5364
rect 4445 5337 4483 5343
rect 4536 5337 4572 5343
rect 4829 5337 4844 5343
rect 4877 5337 4892 5343
rect 5464 5336 5468 5344
rect 5532 5343 5540 5344
rect 5532 5337 5548 5343
rect 1197 5317 1235 5323
rect 1277 5317 1308 5323
rect 1325 5317 1379 5323
rect 1389 5317 1420 5323
rect 1453 5317 1484 5323
rect 1677 5317 1692 5323
rect 2564 5317 2643 5323
rect 3636 5317 3667 5323
rect 3684 5317 3708 5323
rect 3748 5317 3763 5323
rect 4301 5323 4307 5336
rect 4253 5317 4307 5323
rect 205 5297 243 5303
rect 1252 5297 1267 5303
rect 1476 5297 1491 5303
rect 1604 5297 1635 5303
rect 2116 5297 2131 5303
rect 3480 5296 3484 5304
rect 4253 5297 4259 5317
rect 4388 5317 4403 5323
rect 4836 5317 4851 5323
rect 4980 5317 4995 5323
rect 5213 5317 5228 5323
rect 5236 5317 5251 5323
rect 5853 5317 5875 5323
rect 5933 5317 5948 5323
rect 5853 5304 5859 5317
rect 4628 5297 4675 5303
rect 5620 5297 5635 5303
rect 228 5277 243 5283
rect 1501 5277 1516 5283
rect 1901 5277 1916 5283
rect 5789 5277 5820 5283
rect 5789 5257 5795 5277
rect 3188 5236 3190 5244
rect 4996 5236 4998 5244
rect 5252 5236 5254 5244
rect 1560 5206 1566 5214
rect 1574 5206 1580 5214
rect 1588 5206 1594 5214
rect 1602 5206 1608 5214
rect 4632 5206 4638 5214
rect 4646 5206 4652 5214
rect 4660 5206 4666 5214
rect 4674 5206 4680 5214
rect 250 5176 252 5184
rect 644 5176 648 5184
rect 1380 5176 1382 5184
rect 1994 5176 1996 5184
rect 2500 5176 2502 5184
rect 3962 5176 3964 5184
rect 5348 5176 5352 5184
rect 6008 5176 6012 5184
rect 909 5137 924 5143
rect 4308 5136 4310 5144
rect 45 5103 51 5123
rect 813 5117 835 5123
rect 964 5116 972 5124
rect 45 5097 60 5103
rect 168 5097 220 5103
rect 388 5097 403 5103
rect 500 5097 515 5103
rect 836 5097 851 5103
rect 1005 5103 1011 5123
rect 973 5097 1011 5103
rect 1037 5097 1052 5103
rect 1188 5097 1219 5103
rect 1405 5103 1411 5123
rect 1901 5117 1916 5123
rect 1956 5117 1971 5123
rect 2148 5117 2163 5123
rect 4045 5117 4060 5123
rect 4413 5117 4428 5123
rect 5636 5117 5651 5123
rect 1405 5097 1420 5103
rect 1428 5097 1443 5103
rect 1933 5097 1964 5103
rect 2196 5097 2227 5103
rect 2452 5097 2499 5103
rect 2813 5097 2828 5103
rect 3229 5097 3260 5103
rect 3405 5097 3420 5103
rect 93 5077 115 5083
rect 93 5064 99 5077
rect 500 5077 531 5083
rect 877 5077 892 5083
rect 1469 5077 1491 5083
rect 1732 5077 1779 5083
rect 2013 5077 2060 5083
rect 2100 5077 2115 5083
rect 2333 5077 2364 5083
rect 2429 5077 2444 5083
rect 2461 5077 2483 5083
rect 493 5057 508 5063
rect 1661 5057 1699 5063
rect 2461 5063 2467 5077
rect 2804 5077 2851 5083
rect 2893 5077 2931 5083
rect 2445 5057 2467 5063
rect 2877 5057 2899 5063
rect 2925 5057 2931 5077
rect 2980 5077 3011 5083
rect 3252 5077 3283 5083
rect 3320 5077 3340 5083
rect 3405 5077 3411 5097
rect 3981 5097 4019 5103
rect 3981 5084 3987 5097
rect 4125 5097 4156 5103
rect 5917 5097 5980 5103
rect 3572 5077 3603 5083
rect 3613 5077 3644 5083
rect 3805 5077 3820 5083
rect 5165 5077 5187 5083
rect 5245 5077 5315 5083
rect 5876 5077 5891 5083
rect 3380 5056 3388 5064
rect 580 5036 582 5044
rect 1524 5036 1528 5044
rect 5128 5036 5132 5044
rect 6132 5036 6136 5044
rect 3112 5006 3118 5014
rect 3126 5006 3132 5014
rect 3140 5006 3146 5014
rect 3154 5006 3160 5014
rect 548 4976 550 4984
rect 612 4976 616 4984
rect 954 4976 956 4984
rect 1533 4977 1596 4983
rect 1666 4977 1708 4983
rect 3112 4976 3116 4984
rect 3316 4976 3320 4984
rect 3540 4977 3555 4983
rect 3860 4976 3862 4984
rect 4186 4976 4188 4984
rect 4714 4976 4716 4984
rect 5188 4976 5190 4984
rect 5524 4976 5526 4984
rect 5565 4977 5580 4983
rect 5789 4977 5804 4983
rect 5988 4977 6003 4983
rect 6052 4976 6054 4984
rect 6116 4976 6120 4984
rect 420 4957 435 4963
rect 1181 4957 1219 4963
rect 1588 4957 1619 4963
rect 2221 4957 2236 4963
rect 3924 4956 3932 4964
rect 4525 4957 4540 4963
rect 4637 4957 4652 4963
rect 829 4923 835 4943
rect 1229 4937 1244 4943
rect 1556 4937 1635 4943
rect 2365 4937 2380 4943
rect 2765 4937 2780 4943
rect 3149 4937 3180 4943
rect 3400 4936 3404 4944
rect 3752 4937 3788 4943
rect 3892 4937 3916 4943
rect 4644 4937 4723 4943
rect 4749 4943 4755 4963
rect 4765 4957 4780 4963
rect 4740 4937 4755 4943
rect 4781 4937 4803 4943
rect 829 4917 867 4923
rect 1005 4917 1043 4923
rect 1085 4917 1123 4923
rect 1197 4917 1212 4923
rect 1037 4904 1043 4917
rect 1492 4917 1507 4923
rect 1636 4917 1651 4923
rect 1853 4917 1884 4923
rect 1949 4917 1964 4923
rect 2557 4917 2572 4923
rect 2637 4923 2643 4936
rect 4781 4924 4787 4937
rect 5245 4937 5267 4943
rect 5309 4937 5324 4943
rect 5416 4936 5420 4944
rect 2637 4917 2675 4923
rect 2749 4917 2796 4923
rect 3588 4917 3603 4923
rect 4100 4917 4115 4923
rect 4845 4917 4883 4923
rect 5300 4917 5331 4923
rect 5596 4917 5612 4923
rect 5596 4912 5604 4917
rect 5964 4912 5972 4916
rect 877 4897 892 4903
rect 1540 4897 1580 4903
rect 2829 4897 2844 4903
rect 2964 4896 2972 4904
rect 4164 4897 4179 4903
rect 5252 4897 5267 4903
rect 5533 4897 5555 4903
rect 5629 4897 5651 4903
rect 5748 4897 5763 4903
rect 5812 4897 5827 4903
rect 5940 4897 5955 4903
rect 280 4876 284 4884
rect 772 4876 776 4884
rect 2045 4877 2060 4883
rect 2068 4877 2092 4883
rect 3204 4877 3251 4883
rect 3629 4877 3644 4883
rect 4884 4876 4886 4884
rect 5652 4877 5683 4883
rect 5965 4883 5971 4903
rect 5933 4877 5971 4883
rect 5933 4857 5939 4877
rect 1332 4836 1334 4844
rect 1988 4836 1990 4844
rect 2618 4836 2620 4844
rect 2906 4836 2908 4844
rect 1560 4806 1566 4814
rect 1574 4806 1580 4814
rect 1588 4806 1594 4814
rect 1602 4806 1608 4814
rect 4632 4806 4638 4814
rect 4646 4806 4652 4814
rect 4660 4806 4666 4814
rect 4674 4806 4680 4814
rect 72 4776 76 4784
rect 740 4776 748 4784
rect 3508 4776 3510 4784
rect 3572 4776 3574 4784
rect 5156 4776 5160 4784
rect 6138 4776 6140 4784
rect 632 4736 636 4744
rect 948 4736 950 4744
rect 1012 4737 1043 4743
rect 1524 4737 1555 4743
rect 1780 4736 1782 4744
rect 2020 4737 2044 4743
rect 2445 4737 2460 4743
rect 3844 4737 3875 4743
rect 5252 4736 5254 4744
rect 1277 4717 1292 4723
rect 2004 4717 2019 4723
rect 3869 4717 3907 4723
rect 4941 4717 4963 4723
rect 4973 4717 5011 4723
rect 5405 4717 5427 4723
rect 5869 4717 5891 4723
rect 5908 4717 5923 4723
rect 340 4697 392 4703
rect 541 4697 579 4703
rect 861 4697 940 4703
rect 189 4683 195 4696
rect 173 4677 195 4683
rect 221 4677 236 4683
rect 196 4657 211 4663
rect 221 4657 227 4677
rect 333 4677 339 4696
rect 573 4677 579 4697
rect 980 4697 995 4703
rect 1172 4697 1251 4703
rect 1565 4697 1644 4703
rect 2925 4697 2956 4703
rect 3940 4697 3987 4703
rect 3997 4697 4012 4703
rect 4076 4703 4084 4708
rect 4076 4697 4099 4703
rect 4157 4697 4179 4703
rect 4173 4684 4179 4697
rect 4420 4697 4435 4703
rect 4445 4697 4476 4703
rect 4669 4697 4739 4703
rect 4733 4684 4739 4697
rect 5405 4697 5420 4703
rect 5613 4697 5635 4703
rect 5725 4697 5756 4703
rect 6164 4697 6179 4703
rect 877 4677 892 4683
rect 909 4677 931 4683
rect 1181 4677 1196 4683
rect 909 4663 915 4677
rect 1204 4677 1235 4683
rect 1432 4677 1475 4683
rect 2120 4677 2140 4683
rect 2349 4677 2364 4683
rect 3108 4677 3171 4683
rect 3293 4677 3324 4683
rect 3389 4677 3404 4683
rect 3956 4677 3971 4683
rect 4189 4677 4204 4683
rect 5341 4677 5356 4683
rect 5453 4677 5484 4683
rect 5597 4677 5612 4683
rect 6077 4677 6092 4683
rect 893 4657 915 4663
rect 1172 4657 1187 4663
rect 2196 4656 2204 4664
rect 2365 4657 2403 4663
rect 3316 4657 3331 4663
rect 3341 4657 3363 4663
rect 3821 4657 3836 4663
rect 276 4636 280 4644
rect 2308 4636 2318 4644
rect 2445 4637 2460 4643
rect 2701 4637 2716 4643
rect 2900 4636 2910 4644
rect 5018 4636 5020 4644
rect 3112 4606 3118 4614
rect 3126 4606 3132 4614
rect 3140 4606 3146 4614
rect 3154 4606 3160 4614
rect 72 4576 76 4584
rect 344 4576 348 4584
rect 824 4576 828 4584
rect 1096 4576 1100 4584
rect 1514 4576 1516 4584
rect 2306 4577 2332 4583
rect 3620 4577 3635 4583
rect 3962 4576 3964 4584
rect 4180 4577 4195 4583
rect 4378 4576 4380 4584
rect 4740 4576 4742 4584
rect 4890 4576 4892 4584
rect 5066 4576 5068 4584
rect 5172 4576 5176 4584
rect 5588 4576 5590 4584
rect 5898 4576 5900 4584
rect 6029 4577 6051 4583
rect 1341 4557 1363 4563
rect 173 4537 195 4543
rect 381 4537 396 4543
rect 1156 4537 1187 4543
rect 765 4523 771 4536
rect 733 4517 771 4523
rect 1181 4517 1187 4537
rect 1213 4537 1260 4543
rect 1325 4537 1340 4543
rect 1357 4543 1363 4557
rect 1757 4557 1779 4563
rect 1357 4537 1379 4543
rect 1741 4537 1756 4543
rect 1773 4543 1779 4557
rect 2244 4557 2259 4563
rect 1773 4537 1795 4543
rect 1309 4517 1324 4523
rect 1332 4517 1395 4523
rect 1645 4517 1660 4523
rect 1732 4517 1811 4523
rect 1837 4517 1875 4523
rect 1901 4517 1916 4523
rect 1837 4504 1843 4517
rect 1876 4496 1884 4504
rect 1901 4497 1907 4517
rect 2205 4517 2268 4523
rect 2413 4523 2419 4543
rect 2740 4537 2755 4543
rect 2765 4537 2780 4543
rect 2925 4543 2931 4563
rect 4429 4557 4451 4563
rect 2893 4537 2931 4543
rect 3748 4537 3795 4543
rect 4036 4537 4051 4543
rect 4061 4537 4092 4543
rect 4264 4537 4284 4543
rect 4381 4537 4396 4543
rect 4653 4537 4700 4543
rect 4813 4537 4828 4543
rect 4957 4537 4995 4543
rect 5012 4537 5043 4543
rect 5284 4537 5299 4543
rect 2413 4517 2444 4523
rect 3037 4517 3052 4523
rect 3732 4517 3811 4523
rect 4317 4523 4323 4536
rect 5469 4543 5475 4563
rect 6045 4563 6051 4577
rect 6045 4557 6067 4563
rect 5437 4537 5475 4543
rect 5485 4537 5507 4543
rect 5645 4537 5667 4543
rect 5773 4537 5804 4543
rect 5853 4537 5884 4543
rect 4317 4517 4339 4523
rect 4397 4517 4412 4523
rect 4637 4517 4716 4523
rect 4804 4517 4835 4523
rect 2356 4497 2371 4503
rect 2452 4496 2460 4504
rect 3837 4497 3859 4503
rect 4829 4497 4835 4517
rect 5389 4517 5420 4523
rect 5565 4523 5571 4536
rect 6120 4537 6172 4543
rect 5549 4517 5571 4523
rect 5796 4517 5811 4523
rect 4893 4497 4931 4503
rect 5604 4497 5619 4503
rect 936 4476 940 4484
rect 1812 4476 1814 4484
rect 1988 4477 2019 4483
rect 3405 4477 3420 4483
rect 3405 4457 3411 4477
rect 682 4436 684 4444
rect 2394 4436 2396 4444
rect 1560 4406 1566 4414
rect 1574 4406 1580 4414
rect 1588 4406 1594 4414
rect 1602 4406 1608 4414
rect 4632 4406 4638 4414
rect 4646 4406 4652 4414
rect 4660 4406 4666 4414
rect 4674 4406 4680 4414
rect 634 4376 636 4384
rect 1012 4376 1014 4384
rect 2756 4376 2758 4384
rect 4532 4376 4536 4384
rect 4772 4376 4776 4384
rect 5384 4376 5388 4384
rect 5498 4376 5500 4384
rect 413 4337 444 4343
rect 2516 4337 2531 4343
rect 2941 4337 2972 4343
rect 3828 4337 3859 4343
rect 5994 4336 5996 4344
rect 228 4317 259 4323
rect 1876 4317 1891 4323
rect 925 4297 1004 4303
rect 1748 4297 1779 4303
rect 2301 4303 2307 4323
rect 3069 4317 3084 4323
rect 3261 4317 3276 4323
rect 3741 4317 3763 4323
rect 4141 4317 4163 4323
rect 4237 4317 4252 4323
rect 2301 4297 2323 4303
rect 29 4277 44 4283
rect 100 4277 131 4283
rect 285 4277 316 4283
rect 516 4277 531 4283
rect 765 4277 780 4283
rect 941 4277 956 4283
rect 973 4277 995 4283
rect 1085 4277 1107 4283
rect 509 4257 531 4263
rect 973 4263 979 4277
rect 1101 4264 1107 4277
rect 1469 4277 1507 4283
rect 2317 4284 2323 4297
rect 2861 4297 2892 4303
rect 3580 4303 3588 4308
rect 3580 4297 3603 4303
rect 3901 4297 3932 4303
rect 4301 4303 4307 4323
rect 4884 4317 4899 4323
rect 5437 4317 5475 4323
rect 5956 4317 5971 4323
rect 4269 4297 4307 4303
rect 4372 4297 4403 4303
rect 4413 4297 4467 4303
rect 6020 4297 6035 4303
rect 6100 4297 6131 4303
rect 1948 4277 1964 4283
rect 1948 4276 1956 4277
rect 2493 4277 2531 4283
rect 957 4257 979 4263
rect 2493 4257 2499 4277
rect 3645 4277 3667 4283
rect 3709 4277 3724 4283
rect 3645 4264 3651 4277
rect 3972 4277 3987 4283
rect 4308 4277 4323 4283
rect 4333 4277 4355 4283
rect 4621 4277 4691 4283
rect 4829 4277 4867 4283
rect 5533 4277 5571 4283
rect 5581 4277 5612 4283
rect 5668 4277 5699 4283
rect 6013 4277 6035 4283
rect 6093 4277 6108 4283
rect 2893 4257 2908 4263
rect 3485 4257 3507 4263
rect 4365 4257 4387 4263
rect 4852 4256 4860 4264
rect 6109 4257 6115 4276
rect 330 4236 332 4244
rect 1066 4236 1068 4244
rect 2077 4237 2092 4243
rect 5172 4236 5176 4244
rect 5780 4236 5784 4244
rect 6196 4236 6200 4244
rect 3112 4206 3118 4214
rect 3126 4206 3132 4214
rect 3140 4206 3146 4214
rect 3154 4206 3160 4214
rect 72 4176 76 4184
rect 184 4176 188 4184
rect 250 4176 252 4184
rect 456 4176 460 4184
rect 994 4176 1004 4184
rect 1028 4177 1059 4183
rect 1508 4176 1510 4184
rect 1748 4176 1752 4184
rect 2820 4177 2835 4183
rect 3373 4177 3388 4183
rect 3844 4176 3846 4184
rect 4554 4176 4556 4184
rect 4632 4177 4684 4183
rect 5389 4177 5404 4183
rect 5949 4177 5964 4183
rect 909 4157 924 4163
rect 1396 4156 1404 4164
rect 1924 4157 1939 4163
rect 2141 4157 2163 4163
rect 5044 4157 5068 4163
rect 5140 4156 5148 4164
rect 596 4137 636 4143
rect 1181 4137 1212 4143
rect 1341 4137 1356 4143
rect 1469 4137 1491 4143
rect 2141 4137 2156 4143
rect 2189 4137 2204 4143
rect 2564 4137 2611 4143
rect 3197 4137 3228 4143
rect 3444 4137 3475 4143
rect 3572 4137 3587 4143
rect 317 4117 332 4123
rect 573 4117 588 4123
rect 596 4117 659 4123
rect 717 4117 732 4123
rect 1309 4117 1324 4123
rect 2029 4117 2076 4123
rect 2317 4117 2355 4123
rect 2548 4117 2627 4123
rect 2765 4117 2780 4123
rect 2925 4117 2940 4123
rect 3220 4117 3235 4123
rect 3501 4117 3516 4123
rect 1517 4097 1539 4103
rect 2669 4097 2684 4103
rect 2900 4097 2915 4103
rect 3213 4097 3219 4116
rect 3453 4097 3468 4103
rect 3501 4097 3507 4117
rect 3965 4123 3971 4143
rect 4788 4137 4803 4143
rect 5085 4137 5107 4143
rect 5101 4124 5107 4137
rect 5149 4137 5164 4143
rect 5549 4143 5555 4163
rect 5764 4157 5779 4163
rect 5517 4137 5555 4143
rect 5565 4137 5587 4143
rect 6052 4137 6067 4143
rect 3940 4117 3971 4123
rect 4765 4117 4780 4123
rect 4788 4117 4819 4123
rect 5037 4117 5052 4123
rect 5252 4117 5267 4123
rect 6036 4117 6083 4123
rect 6116 4117 6147 4123
rect 6180 4117 6195 4123
rect 3693 4097 3708 4103
rect 4717 4097 4739 4103
rect 4756 4096 4764 4104
rect 5428 4097 5443 4103
rect 5981 4097 5996 4103
rect 1516 4084 1524 4088
rect 4676 4077 4723 4083
rect 5412 4077 5475 4083
rect 5789 4077 5843 4083
rect 5853 4077 5884 4083
rect 1844 4036 1846 4044
rect 1908 4036 1910 4044
rect 2756 4036 2758 4044
rect 3117 4037 3164 4043
rect 6026 4036 6028 4044
rect 6084 4036 6086 4044
rect 6196 4036 6198 4044
rect 1560 4006 1566 4014
rect 1574 4006 1580 4014
rect 1588 4006 1594 4014
rect 1602 4006 1608 4014
rect 4632 4006 4638 4014
rect 4646 4006 4652 4014
rect 4660 4006 4666 4014
rect 4674 4006 4680 4014
rect 72 3976 76 3984
rect 452 3976 454 3984
rect 794 3976 796 3984
rect 852 3976 854 3984
rect 916 3976 918 3984
rect 1098 3976 1100 3984
rect 1204 3976 1206 3984
rect 1332 3976 1334 3984
rect 2650 3976 2652 3984
rect 3085 3977 3132 3983
rect 3284 3976 3286 3984
rect 3348 3976 3350 3984
rect 4776 3976 4780 3984
rect 5610 3976 5612 3984
rect 980 3936 982 3944
rect 2330 3936 2332 3944
rect 2748 3937 2764 3943
rect 2748 3932 2756 3937
rect 3021 3937 3075 3943
rect 3924 3936 3926 3944
rect 4052 3937 4131 3943
rect 4845 3937 4860 3943
rect 5748 3937 5763 3943
rect 5892 3937 5923 3943
rect 3068 3924 3076 3928
rect 349 3917 371 3923
rect 477 3917 499 3923
rect 516 3917 531 3923
rect 733 3917 771 3923
rect 1005 3917 1043 3923
rect 372 3897 387 3903
rect 420 3897 451 3903
rect 484 3897 499 3903
rect 813 3897 851 3903
rect 813 3884 819 3897
rect 925 3897 956 3903
rect 1229 3903 1235 3923
rect 1357 3917 1395 3923
rect 1405 3917 1420 3923
rect 1229 3897 1267 3903
rect 1501 3897 1523 3903
rect 1565 3897 1612 3903
rect 2052 3897 2131 3903
rect 2141 3897 2156 3903
rect 2333 3897 2371 3903
rect 2861 3903 2867 3923
rect 2989 3917 3004 3923
rect 3540 3916 3548 3924
rect 2861 3897 2876 3903
rect 3108 3897 3171 3903
rect 3181 3897 3196 3903
rect 3869 3897 3900 3903
rect 4621 3903 4627 3923
rect 4925 3917 4947 3923
rect 5197 3917 5212 3923
rect 5252 3917 5267 3923
rect 5668 3916 5676 3924
rect 5917 3917 5955 3923
rect 6061 3917 6067 3936
rect 4596 3897 4627 3903
rect 5085 3897 5100 3903
rect 5204 3897 5235 3903
rect 5332 3897 5347 3903
rect 5405 3897 5427 3903
rect 5421 3884 5427 3897
rect 6189 3897 6220 3903
rect 292 3877 323 3883
rect 420 3877 435 3883
rect 605 3877 636 3883
rect 1149 3877 1187 3883
rect 1300 3877 1315 3883
rect 1524 3877 1539 3883
rect 1565 3877 1651 3883
rect 292 3857 307 3863
rect 1565 3857 1571 3877
rect 1837 3877 1884 3883
rect 2068 3877 2115 3883
rect 3252 3877 3267 3883
rect 3805 3877 3836 3883
rect 4813 3877 4828 3883
rect 5716 3877 5731 3883
rect 6084 3877 6099 3883
rect 6205 3877 6236 3883
rect 1645 3857 1683 3863
rect 1768 3836 1772 3844
rect 2456 3836 2460 3844
rect 4634 3836 4636 3844
rect 5805 3837 5820 3843
rect 5869 3837 5884 3843
rect 5972 3837 5987 3843
rect 6029 3837 6044 3843
rect 3112 3806 3118 3814
rect 3126 3806 3132 3814
rect 3140 3806 3146 3814
rect 3154 3806 3160 3814
rect 52 3776 56 3784
rect 212 3776 214 3784
rect 538 3776 540 3784
rect 1581 3777 1628 3783
rect 2634 3776 2636 3784
rect 2788 3776 2790 3784
rect 3514 3776 3516 3784
rect 3896 3776 3900 3784
rect 4436 3776 4438 3784
rect 4506 3776 4508 3784
rect 5320 3776 5324 3784
rect 644 3756 652 3764
rect 1005 3757 1020 3763
rect 109 3737 140 3743
rect 484 3737 499 3743
rect 717 3737 732 3743
rect 925 3737 956 3743
rect 1069 3743 1075 3763
rect 2516 3757 2531 3763
rect 1037 3737 1075 3743
rect 1172 3737 1187 3743
rect 445 3717 476 3723
rect 637 3717 675 3723
rect 701 3717 716 3723
rect 669 3697 675 3717
rect 852 3717 867 3723
rect 964 3717 979 3723
rect 1325 3723 1331 3743
rect 2669 3743 2675 3763
rect 2685 3757 2707 3763
rect 2660 3737 2675 3743
rect 2909 3737 2924 3743
rect 2989 3737 3004 3743
rect 3229 3743 3235 3763
rect 3373 3757 3404 3763
rect 3661 3757 3699 3763
rect 3197 3737 3235 3743
rect 3268 3737 3292 3743
rect 3325 3737 3340 3743
rect 3988 3737 4003 3743
rect 4340 3737 4355 3743
rect 4525 3737 4547 3743
rect 4653 3737 4723 3743
rect 4733 3737 4771 3743
rect 4717 3724 4723 3737
rect 4877 3737 4908 3743
rect 4948 3737 4963 3743
rect 5037 3737 5084 3743
rect 5181 3737 5203 3743
rect 5789 3743 5795 3763
rect 5716 3737 5731 3743
rect 5789 3737 5804 3743
rect 5997 3737 6012 3743
rect 6088 3737 6108 3743
rect 6164 3737 6179 3743
rect 6205 3737 6220 3743
rect 1261 3717 1331 3723
rect 1380 3717 1395 3723
rect 1405 3717 1443 3723
rect 1389 3704 1395 3717
rect 1437 3704 1443 3717
rect 1517 3717 1548 3723
rect 1917 3717 1948 3723
rect 2077 3717 2092 3723
rect 2429 3717 2467 3723
rect 3309 3717 3347 3723
rect 3540 3717 3555 3723
rect 3965 3717 3996 3723
rect 1588 3697 1628 3703
rect 2045 3697 2083 3703
rect 2173 3697 2188 3703
rect 2797 3697 2819 3703
rect 3092 3696 3100 3704
rect 4813 3697 4835 3703
rect 4989 3697 5004 3703
rect 5677 3697 5699 3703
rect 6029 3697 6051 3703
rect 2461 3677 2492 3683
rect 1178 3636 1180 3644
rect 1272 3636 1276 3644
rect 1704 3636 1708 3644
rect 3194 3636 3196 3644
rect 1560 3606 1566 3614
rect 1574 3606 1580 3614
rect 1588 3606 1594 3614
rect 1602 3606 1608 3614
rect 4632 3606 4638 3614
rect 4646 3606 4652 3614
rect 4660 3606 4666 3614
rect 4674 3606 4680 3614
rect 72 3576 76 3584
rect 180 3576 182 3584
rect 308 3576 310 3584
rect 362 3576 364 3584
rect 564 3576 566 3584
rect 804 3576 806 3584
rect 2052 3576 2054 3584
rect 2436 3576 2438 3584
rect 2660 3576 2662 3584
rect 3476 3576 3478 3584
rect 3834 3576 3836 3584
rect 3960 3576 3964 3584
rect 4202 3576 4204 3584
rect 4612 3576 4616 3584
rect 5114 3576 5116 3584
rect 5172 3576 5174 3584
rect 5434 3576 5436 3584
rect 6004 3576 6008 3584
rect 5514 3556 5516 3564
rect 458 3536 460 3544
rect 1341 3537 1356 3543
rect 1380 3537 1395 3543
rect 1620 3536 1622 3544
rect 1796 3537 1827 3543
rect 2356 3537 2387 3543
rect 4308 3536 4310 3544
rect 5732 3537 5747 3543
rect 6196 3537 6211 3543
rect 205 3503 211 3523
rect 1220 3517 1235 3523
rect 1940 3514 1944 3522
rect 2548 3516 2556 3524
rect 205 3497 243 3503
rect 253 3497 268 3503
rect 276 3497 307 3503
rect 340 3497 355 3503
rect 484 3497 499 3503
rect 724 3497 739 3503
rect 749 3497 780 3503
rect 836 3497 851 3503
rect 1044 3497 1116 3503
rect 1405 3497 1420 3503
rect 1533 3497 1596 3503
rect 477 3477 492 3483
rect 637 3477 675 3483
rect 701 3477 723 3483
rect 701 3464 707 3477
rect 1060 3477 1107 3483
rect 1572 3477 1603 3483
rect 1725 3483 1731 3503
rect 1837 3497 1852 3503
rect 1981 3497 2044 3503
rect 1981 3484 1987 3497
rect 2084 3497 2115 3503
rect 2397 3497 2412 3503
rect 2573 3503 2579 3523
rect 2532 3497 2547 3503
rect 2573 3497 2659 3503
rect 3300 3497 3315 3503
rect 3396 3497 3411 3503
rect 3501 3503 3507 3523
rect 3789 3517 3811 3523
rect 4066 3516 4076 3524
rect 4164 3517 4179 3523
rect 4749 3517 4764 3523
rect 5252 3517 5267 3523
rect 3501 3497 3539 3503
rect 3652 3497 3676 3503
rect 3837 3497 3891 3503
rect 4797 3497 4835 3503
rect 5133 3497 5164 3503
rect 1700 3477 1731 3483
rect 1757 3477 1772 3483
rect 2013 3477 2028 3483
rect 2013 3463 2019 3477
rect 2788 3477 2804 3483
rect 2796 3476 2804 3477
rect 4004 3477 4019 3483
rect 4141 3477 4156 3483
rect 4669 3477 4700 3483
rect 4852 3477 4867 3483
rect 5005 3477 5027 3483
rect 5133 3477 5139 3497
rect 5245 3484 5251 3503
rect 5485 3497 5500 3503
rect 5645 3503 5651 3523
rect 5700 3517 5715 3523
rect 5908 3517 5923 3523
rect 5540 3497 5571 3503
rect 5645 3497 5683 3503
rect 6068 3497 6083 3503
rect 5533 3477 5555 3483
rect 5597 3477 5619 3483
rect 5533 3464 5539 3477
rect 5956 3477 5971 3483
rect 6077 3477 6083 3497
rect 6148 3497 6179 3503
rect 6173 3477 6179 3497
rect 6205 3477 6220 3483
rect 1972 3457 1987 3463
rect 1997 3457 2019 3463
rect 4692 3457 4739 3463
rect 1012 3436 1022 3444
rect 2868 3436 2872 3444
rect 3028 3437 3043 3443
rect 3140 3437 3187 3443
rect 6116 3436 6120 3444
rect 3112 3406 3118 3414
rect 3126 3406 3132 3414
rect 3140 3406 3146 3414
rect 3154 3406 3160 3414
rect 186 3376 188 3384
rect 234 3376 236 3384
rect 1512 3376 1516 3384
rect 2349 3377 2364 3383
rect 2957 3377 2972 3383
rect 3274 3376 3276 3384
rect 4324 3376 4328 3384
rect 4458 3376 4460 3384
rect 4792 3376 4796 3384
rect 4996 3376 4998 3384
rect 5044 3376 5046 3384
rect 6068 3376 6072 3384
rect 29 3337 67 3343
rect 228 3337 243 3343
rect 765 3343 771 3363
rect 765 3337 780 3343
rect 893 3337 931 3343
rect 1133 3343 1139 3363
rect 1364 3356 1372 3364
rect 2861 3357 2883 3363
rect 3181 3357 3196 3363
rect 3332 3357 3347 3363
rect 4068 3357 4092 3363
rect 1101 3337 1139 3343
rect 1165 3337 1219 3343
rect 1629 3337 1644 3343
rect 1876 3337 1891 3343
rect 2260 3337 2275 3343
rect 3348 3337 3363 3343
rect 612 3317 627 3323
rect 637 3317 675 3323
rect 973 3317 1011 3323
rect 1021 3317 1075 3323
rect 973 3297 979 3317
rect 1709 3317 1740 3323
rect 1901 3317 1916 3323
rect 2237 3317 2284 3323
rect 3085 3317 3148 3323
rect 3245 3317 3260 3323
rect 3597 3323 3603 3343
rect 3636 3337 3651 3343
rect 3580 3317 3603 3323
rect 3580 3312 3588 3317
rect 3901 3317 3923 3323
rect 4125 3323 4131 3343
rect 4285 3323 4291 3343
rect 4525 3343 4531 3363
rect 4637 3357 4707 3363
rect 4941 3344 4947 3363
rect 5108 3357 5139 3363
rect 4477 3337 4499 3343
rect 4525 3337 4540 3343
rect 4493 3324 4499 3337
rect 4589 3337 4604 3343
rect 4909 3337 4940 3343
rect 5012 3337 5027 3343
rect 5261 3343 5267 3356
rect 5060 3337 5091 3343
rect 5133 3337 5171 3343
rect 5261 3337 5283 3343
rect 4116 3317 4131 3323
rect 4253 3317 4291 3323
rect 4413 3317 4451 3323
rect 1837 3297 1884 3303
rect 1917 3297 1932 3303
rect 2029 3297 2044 3303
rect 2141 3297 2156 3303
rect 3517 3297 3539 3303
rect 3629 3297 3644 3303
rect 4445 3297 4451 3317
rect 4573 3317 4611 3323
rect 5460 3317 5491 3323
rect 5837 3323 5843 3363
rect 5821 3317 5843 3323
rect 5821 3304 5827 3317
rect 5949 3317 5980 3323
rect 6029 3323 6035 3343
rect 6173 3337 6211 3343
rect 5997 3317 6035 3323
rect 6173 3317 6179 3337
rect 5005 3297 5020 3303
rect 5389 3297 5411 3303
rect 5565 3297 5580 3303
rect 1018 3276 1020 3284
rect 1060 3277 1075 3283
rect 1812 3276 1814 3284
rect 4957 3277 4972 3283
rect 3085 3257 3132 3263
rect 1748 3236 1750 3244
rect 2004 3236 2006 3244
rect 2746 3236 2748 3244
rect 4184 3236 4188 3244
rect 5242 3236 5244 3244
rect 6164 3236 6166 3244
rect 1560 3206 1566 3214
rect 1574 3206 1580 3214
rect 1588 3206 1594 3214
rect 1602 3206 1608 3214
rect 4632 3206 4638 3214
rect 4646 3206 4652 3214
rect 4660 3206 4666 3214
rect 4674 3206 4680 3214
rect 394 3176 396 3184
rect 564 3176 566 3184
rect 900 3176 902 3184
rect 1188 3176 1190 3184
rect 1812 3176 1814 3184
rect 2260 3176 2262 3184
rect 2938 3176 2940 3184
rect 3162 3176 3164 3184
rect 3220 3176 3222 3184
rect 3716 3176 3718 3184
rect 4570 3176 4572 3184
rect 4858 3176 4860 3184
rect 4932 3176 4936 3184
rect 5268 3176 5270 3184
rect 5476 3176 5478 3184
rect 5844 3176 5846 3184
rect 5914 3176 5916 3184
rect 5972 3176 5974 3184
rect 836 3136 838 3144
rect 1836 3137 1891 3143
rect 2061 3137 2092 3143
rect 2653 3143 2659 3163
rect 2653 3137 2723 3143
rect 3300 3137 3331 3143
rect 3405 3137 3420 3143
rect 3540 3136 3542 3144
rect 3604 3137 3619 3143
rect 3796 3137 3811 3143
rect 4100 3137 4115 3143
rect 5380 3136 5384 3144
rect 5725 3137 5779 3143
rect 364 3132 372 3136
rect 2716 3124 2724 3128
rect 5724 3124 5732 3128
rect 212 3117 227 3123
rect 676 3114 680 3122
rect 2029 3117 2044 3123
rect 2125 3117 2140 3123
rect 2493 3117 2515 3123
rect 3284 3117 3299 3123
rect 420 3097 435 3103
rect 109 3077 147 3083
rect 260 3077 275 3083
rect 461 3077 476 3083
rect 180 3056 188 3064
rect 356 3057 380 3063
rect 461 3057 467 3077
rect 605 3077 652 3083
rect 957 3077 972 3083
rect 1021 3083 1027 3103
rect 2205 3097 2259 3103
rect 2957 3097 2995 3103
rect 1021 3077 1052 3083
rect 1437 3077 1452 3083
rect 1996 3077 2012 3083
rect 1996 3076 2004 3077
rect 2413 3077 2444 3083
rect 2548 3077 2563 3083
rect 2349 3057 2371 3063
rect 2557 3057 2563 3077
rect 2957 3077 2963 3097
rect 3165 3097 3212 3103
rect 3741 3103 3747 3123
rect 4285 3117 4307 3123
rect 3661 3097 3715 3103
rect 3741 3097 3779 3103
rect 4333 3097 4412 3103
rect 4541 3103 4547 3123
rect 5549 3117 5587 3123
rect 4509 3097 4547 3103
rect 4596 3097 4627 3103
rect 4813 3097 4828 3103
rect 5060 3097 5075 3103
rect 5085 3097 5107 3103
rect 5277 3097 5315 3103
rect 5812 3097 5843 3103
rect 5917 3097 5964 3103
rect 3181 3077 3196 3083
rect 3908 3077 3939 3083
rect 4356 3077 4403 3083
rect 5188 3077 5203 3083
rect 2765 3057 2787 3063
rect 3405 3057 3420 3063
rect 4260 3057 4275 3063
rect 4756 3056 4764 3064
rect 5021 3057 5059 3063
rect 5117 3057 5139 3063
rect 5197 3057 5203 3077
rect 5933 3077 5948 3083
rect 5213 3057 5251 3063
rect 2164 3036 2166 3044
rect 2212 3036 2214 3044
rect 2728 3036 2732 3044
rect 3112 3006 3118 3014
rect 3126 3006 3132 3014
rect 3140 3006 3146 3014
rect 3154 3006 3160 3014
rect 100 2976 104 2984
rect 266 2976 268 2984
rect 618 2976 620 2984
rect 858 2976 860 2984
rect 1336 2976 1340 2984
rect 1565 2977 1612 2983
rect 2797 2977 2812 2983
rect 3108 2977 3155 2983
rect 3716 2976 3718 2984
rect 4888 2976 4892 2984
rect 5434 2976 5436 2984
rect 6090 2976 6092 2984
rect 3716 2957 3747 2963
rect 4589 2957 4611 2963
rect 61 2923 67 2943
rect 1261 2937 1283 2943
rect 29 2917 67 2923
rect 877 2917 900 2923
rect 892 2912 900 2917
rect 1076 2917 1107 2923
rect 1261 2923 1267 2937
rect 1588 2937 1635 2943
rect 1768 2937 1788 2943
rect 2196 2937 2211 2943
rect 2637 2937 2652 2943
rect 2916 2937 2947 2943
rect 3748 2937 3763 2943
rect 3860 2937 3891 2943
rect 3965 2937 3987 2943
rect 4184 2936 4188 2944
rect 4356 2937 4371 2943
rect 1236 2917 1267 2923
rect 2180 2917 2227 2923
rect 2237 2917 2268 2923
rect 2628 2917 2675 2923
rect 2828 2917 2851 2923
rect 2828 2912 2836 2917
rect 3373 2917 3404 2923
rect 3453 2917 3484 2923
rect 4308 2917 4323 2923
rect 4333 2917 4380 2923
rect 4445 2917 4460 2923
rect 4829 2923 4835 2943
rect 5197 2943 5203 2963
rect 5485 2957 5507 2963
rect 5748 2956 5756 2964
rect 5885 2957 5900 2963
rect 5197 2937 5267 2943
rect 5357 2924 5363 2943
rect 5933 2943 5939 2956
rect 5933 2937 5955 2943
rect 4797 2917 4835 2923
rect 5156 2917 5187 2923
rect 5364 2917 5395 2923
rect 6045 2917 6060 2923
rect 548 2897 563 2903
rect 1218 2896 1228 2904
rect 1565 2897 1612 2903
rect 3012 2897 3027 2903
rect 3277 2897 3292 2903
rect 3469 2897 3484 2903
rect 3629 2897 3667 2903
rect 3677 2897 3715 2903
rect 3789 2897 3811 2903
rect 3917 2897 3939 2903
rect 4228 2897 4243 2903
rect 4724 2897 4739 2903
rect 5108 2897 5123 2903
rect 412 2884 420 2888
rect 1972 2877 1987 2883
rect 2676 2876 2678 2884
rect 2700 2877 2755 2883
rect 3549 2877 3564 2883
rect 4189 2877 4252 2883
rect 6196 2877 6211 2883
rect 1044 2836 1046 2844
rect 1418 2836 1420 2844
rect 2170 2836 2172 2844
rect 2618 2836 2620 2844
rect 3604 2836 3606 2844
rect 4388 2836 4390 2844
rect 5300 2836 5304 2844
rect 5972 2836 5974 2844
rect 1560 2806 1566 2814
rect 1574 2806 1580 2814
rect 1588 2806 1594 2814
rect 1602 2806 1608 2814
rect 4632 2806 4638 2814
rect 4646 2806 4652 2814
rect 4660 2806 4666 2814
rect 4674 2806 4680 2814
rect 2746 2776 2748 2784
rect 2852 2776 2854 2784
rect 900 2737 931 2743
rect 3204 2737 3219 2743
rect 3933 2737 3964 2743
rect 4436 2736 4438 2744
rect 4516 2737 4547 2743
rect 1661 2717 1676 2723
rect 2573 2717 2588 2723
rect 2996 2717 3011 2723
rect 3028 2717 3043 2723
rect 3108 2717 3123 2723
rect 349 2697 364 2703
rect 660 2697 684 2703
rect 877 2697 908 2703
rect 1037 2697 1052 2703
rect 292 2677 307 2683
rect 1037 2677 1043 2697
rect 1700 2697 1715 2703
rect 2509 2697 2547 2703
rect 2557 2697 2572 2703
rect 2765 2697 2780 2703
rect 1236 2677 1251 2683
rect 1773 2677 1811 2683
rect 1892 2677 1923 2683
rect 2045 2677 2060 2683
rect 2248 2676 2252 2684
rect 2280 2676 2284 2684
rect 2765 2677 2771 2697
rect 3405 2703 3411 2723
rect 3428 2716 3436 2724
rect 3565 2717 3587 2723
rect 3645 2717 3699 2723
rect 3901 2717 3939 2723
rect 4541 2717 4547 2737
rect 5204 2737 5244 2743
rect 3373 2697 3411 2703
rect 3437 2697 3468 2703
rect 3476 2697 3491 2703
rect 3629 2697 3644 2703
rect 3709 2697 3740 2703
rect 3757 2697 3772 2703
rect 4252 2703 4260 2708
rect 4252 2697 4275 2703
rect 4708 2697 4723 2703
rect 4877 2703 4883 2723
rect 5021 2717 5036 2723
rect 5229 2717 5283 2723
rect 5556 2716 5564 2724
rect 4845 2697 4883 2703
rect 4893 2697 4931 2703
rect 5053 2697 5068 2703
rect 4925 2684 4931 2697
rect 5325 2697 5340 2703
rect 5468 2703 5476 2708
rect 5380 2697 5395 2703
rect 5453 2697 5476 2703
rect 5805 2697 5820 2703
rect 5908 2697 5939 2703
rect 5997 2697 6012 2703
rect 3453 2677 3468 2683
rect 3581 2677 3619 2683
rect 3732 2677 3747 2683
rect 4116 2677 4147 2683
rect 4621 2677 4707 2683
rect 4733 2677 4748 2683
rect 845 2657 876 2663
rect 1837 2657 1875 2663
rect 2637 2657 2659 2663
rect 4637 2657 4652 2663
rect 4701 2657 4707 2677
rect 5320 2677 5347 2683
rect 5396 2677 5411 2683
rect 5821 2677 5843 2683
rect 5853 2677 5875 2683
rect 5885 2677 5900 2683
rect 5837 2664 5843 2677
rect 6061 2677 6099 2683
rect 122 2636 124 2644
rect 276 2636 278 2644
rect 1018 2636 1020 2644
rect 3258 2636 3260 2644
rect 3306 2636 3308 2644
rect 4788 2636 4790 2644
rect 5434 2636 5436 2644
rect 5492 2637 5507 2643
rect 3112 2606 3118 2614
rect 3126 2606 3132 2614
rect 3140 2606 3146 2614
rect 3154 2606 3160 2614
rect 813 2577 828 2583
rect 1076 2576 1078 2584
rect 1581 2577 1628 2583
rect 2634 2576 2636 2584
rect 3940 2576 3942 2584
rect 4148 2577 4163 2583
rect 4506 2576 4508 2584
rect 1108 2556 1116 2564
rect 356 2537 371 2543
rect 541 2537 556 2543
rect 868 2537 883 2543
rect 980 2537 995 2543
rect 1165 2537 1187 2543
rect 1620 2537 1651 2543
rect 1741 2537 1763 2543
rect 2061 2543 2067 2563
rect 4388 2557 4403 2563
rect 2004 2537 2035 2543
rect 2061 2537 2099 2543
rect 2717 2537 2732 2543
rect 3053 2537 3116 2543
rect 3236 2537 3267 2543
rect 3277 2537 3331 2543
rect 3357 2537 3372 2543
rect 3533 2537 3548 2543
rect 3588 2537 3619 2543
rect 4340 2537 4355 2543
rect 4365 2537 4396 2543
rect 4660 2537 4723 2543
rect 476 2517 499 2523
rect 476 2512 484 2517
rect 909 2517 924 2523
rect 964 2517 1011 2523
rect 1452 2517 1475 2523
rect 1517 2517 1532 2523
rect 1452 2512 1460 2517
rect 1748 2517 1763 2523
rect 1812 2517 1843 2523
rect 2653 2517 2691 2523
rect 2653 2504 2659 2517
rect 2708 2517 2755 2523
rect 3245 2517 3260 2523
rect 3373 2517 3388 2523
rect 3540 2517 3555 2523
rect 1444 2497 1459 2503
rect 2484 2497 2499 2503
rect 2605 2497 2627 2503
rect 2692 2496 2700 2504
rect 2781 2497 2819 2503
rect 2948 2497 2963 2503
rect 3549 2497 3555 2517
rect 3693 2497 3699 2536
rect 4317 2517 4339 2523
rect 4317 2504 4323 2517
rect 4468 2517 4499 2523
rect 4493 2497 4499 2517
rect 4637 2517 4732 2523
rect 4909 2523 4915 2543
rect 5037 2543 5043 2563
rect 5101 2557 5139 2563
rect 5309 2557 5347 2563
rect 5037 2537 5075 2543
rect 5220 2537 5235 2543
rect 5421 2537 5436 2543
rect 5453 2537 5468 2543
rect 5844 2537 5875 2543
rect 6093 2537 6108 2543
rect 4772 2517 4787 2523
rect 4596 2497 4611 2503
rect 1352 2476 1356 2484
rect 2212 2477 2259 2483
rect 1012 2456 1014 2464
rect 2132 2456 2134 2464
rect 2253 2457 2259 2477
rect 2580 2477 2595 2483
rect 2813 2477 2867 2483
rect 3124 2477 3155 2483
rect 3149 2457 3155 2477
rect 4109 2477 4163 2483
rect 4634 2476 4636 2484
rect 4829 2483 4835 2523
rect 4909 2517 4932 2523
rect 4924 2512 4932 2517
rect 5117 2517 5132 2523
rect 5197 2517 5244 2523
rect 6036 2517 6067 2523
rect 6084 2517 6131 2523
rect 5188 2496 5196 2504
rect 5748 2497 5763 2503
rect 5796 2497 5811 2503
rect 6164 2497 6179 2503
rect 4804 2477 4835 2483
rect 5252 2476 5254 2484
rect 5348 2477 5363 2483
rect 5656 2476 5660 2484
rect 954 2436 956 2444
rect 1668 2436 1670 2444
rect 1844 2436 1846 2444
rect 4020 2436 4022 2444
rect 4740 2436 4742 2444
rect 5972 2436 5976 2444
rect 1560 2406 1566 2414
rect 1574 2406 1580 2414
rect 1588 2406 1594 2414
rect 1602 2406 1608 2414
rect 4632 2406 4638 2414
rect 4646 2406 4652 2414
rect 4660 2406 4666 2414
rect 4674 2406 4680 2414
rect 4810 2376 4812 2384
rect 5668 2376 5670 2384
rect 6084 2376 6086 2384
rect 100 2337 116 2343
rect 108 2332 116 2337
rect 660 2336 662 2344
rect 1908 2336 1910 2344
rect 2333 2337 2364 2343
rect 2692 2337 2716 2343
rect 2820 2337 2844 2343
rect 2900 2337 2931 2343
rect 3972 2337 3987 2343
rect 5220 2336 5224 2344
rect 5533 2337 5564 2343
rect 5853 2337 5868 2343
rect 173 2297 188 2303
rect 765 2303 771 2323
rect 836 2316 844 2324
rect 2493 2317 2547 2323
rect 2781 2317 2835 2323
rect 733 2297 771 2303
rect 893 2297 908 2303
rect 1212 2303 1220 2308
rect 1212 2297 1235 2303
rect 1437 2297 1452 2303
rect 1549 2297 1644 2303
rect 1740 2303 1748 2308
rect 1740 2297 1763 2303
rect 1869 2297 1884 2303
rect 2989 2303 2995 2323
rect 3117 2317 3164 2323
rect 3396 2317 3411 2323
rect 3668 2317 3683 2323
rect 3853 2317 3875 2323
rect 3949 2317 3964 2323
rect 2989 2297 3004 2303
rect 3101 2297 3180 2303
rect 3597 2297 3635 2303
rect 3693 2297 3724 2303
rect 93 2277 108 2283
rect 3629 2284 3635 2297
rect 3997 2303 4003 2323
rect 5053 2317 5075 2323
rect 5757 2317 5772 2323
rect 5949 2317 6003 2323
rect 3997 2297 4028 2303
rect 4637 2303 4643 2316
rect 4637 2297 4723 2303
rect 4772 2297 4787 2303
rect 5309 2297 5324 2303
rect 5629 2297 5660 2303
rect 605 2277 643 2283
rect 1076 2277 1107 2283
rect 1428 2277 1459 2283
rect 1572 2277 1635 2283
rect 2221 2277 2252 2283
rect 2396 2277 2412 2283
rect 2396 2276 2404 2277
rect 2996 2277 3027 2283
rect 3140 2277 3187 2283
rect 3229 2277 3244 2283
rect 3524 2277 3555 2283
rect 3709 2277 3763 2283
rect 4445 2277 4483 2283
rect 4525 2277 4563 2283
rect 932 2256 940 2264
rect 1277 2257 1299 2263
rect 2125 2257 2147 2263
rect 4477 2257 4483 2277
rect 4557 2257 4563 2277
rect 4637 2277 4652 2283
rect 4836 2277 4851 2283
rect 5060 2277 5075 2283
rect 5101 2277 5116 2283
rect 5124 2277 5139 2283
rect 5332 2277 5347 2283
rect 5453 2277 5468 2283
rect 6221 2277 6236 2283
rect 5476 2256 5484 2264
rect 5917 2257 5932 2263
rect 26 2236 28 2244
rect 74 2236 76 2244
rect 317 2237 332 2243
rect 474 2236 476 2244
rect 964 2236 968 2244
rect 1341 2237 1356 2243
rect 1709 2237 1724 2243
rect 2026 2236 2028 2244
rect 2872 2236 2876 2244
rect 3546 2236 3548 2244
rect 4276 2237 4291 2243
rect 4394 2236 4396 2244
rect 4904 2236 4908 2244
rect 6164 2236 6168 2244
rect 3112 2206 3118 2214
rect 3126 2206 3132 2214
rect 3140 2206 3146 2214
rect 3154 2206 3160 2214
rect 680 2176 684 2184
rect 2666 2176 2668 2184
rect 2952 2176 2956 2184
rect 2986 2176 2988 2184
rect 4632 2177 4684 2183
rect 5130 2176 5132 2184
rect 5876 2176 5878 2184
rect 925 2157 947 2163
rect 2884 2156 2892 2164
rect 180 2137 195 2143
rect 301 2143 307 2156
rect 301 2137 323 2143
rect 564 2137 579 2143
rect 1165 2137 1203 2143
rect 1444 2137 1459 2143
rect 2461 2137 2499 2143
rect 2541 2137 2572 2143
rect 2692 2137 2707 2143
rect 2852 2137 2867 2143
rect 3716 2137 3731 2143
rect 3757 2143 3763 2163
rect 3748 2137 3763 2143
rect 3789 2137 3811 2143
rect 3789 2124 3795 2137
rect 4749 2143 4755 2163
rect 5181 2157 5203 2163
rect 5805 2157 5827 2163
rect 5837 2144 5843 2163
rect 5924 2157 5955 2163
rect 4717 2137 4755 2143
rect 5133 2137 5148 2143
rect 5597 2137 5628 2143
rect 5844 2137 5859 2143
rect 5892 2137 5907 2143
rect 5965 2137 6003 2143
rect 6104 2137 6124 2143
rect 6173 2137 6204 2143
rect 324 2117 339 2123
rect 388 2117 403 2123
rect 413 2117 428 2123
rect 548 2117 595 2123
rect 893 2117 908 2123
rect 1261 2117 1299 2123
rect 1428 2117 1475 2123
rect 1485 2117 1500 2123
rect 2397 2117 2412 2123
rect 2621 2117 2659 2123
rect 765 2097 780 2103
rect 1741 2097 1795 2103
rect 2276 2097 2291 2103
rect 2653 2097 2659 2117
rect 3012 2117 3027 2123
rect 3885 2117 3900 2123
rect 4365 2117 4396 2123
rect 4676 2117 4700 2123
rect 4925 2117 4940 2123
rect 5357 2117 5388 2123
rect 5740 2117 5763 2123
rect 5740 2112 5748 2117
rect 2740 2097 2755 2103
rect 2845 2097 2883 2103
rect 3684 2097 3699 2103
rect 4765 2097 4787 2103
rect 620 2077 675 2083
rect 772 2077 803 2083
rect 1364 2077 1396 2083
rect 1500 2077 1555 2083
rect 1565 2077 1644 2083
rect 2260 2077 2323 2083
rect 2580 2077 2595 2083
rect 2892 2083 2900 2088
rect 2820 2077 2835 2083
rect 2892 2077 2924 2083
rect 3092 2077 3107 2083
rect 3213 2077 3244 2083
rect 1108 2056 1112 2064
rect 3213 2057 3219 2077
rect 3549 2077 3564 2083
rect 4333 2077 4348 2083
rect 4573 2077 4604 2083
rect 4973 2077 4988 2083
rect 5492 2077 5555 2083
rect 340 2036 342 2044
rect 3117 2037 3164 2043
rect 4922 2036 4924 2044
rect 1560 2006 1566 2014
rect 1574 2006 1580 2014
rect 1588 2006 1594 2014
rect 1602 2006 1608 2014
rect 4632 2006 4638 2014
rect 4646 2006 4652 2014
rect 4660 2006 4666 2014
rect 4674 2006 4680 2014
rect 980 1976 982 1984
rect 1300 1976 1302 1984
rect 3434 1976 3436 1984
rect 3626 1976 3628 1984
rect 253 1937 268 1943
rect 1236 1937 1251 1943
rect 2429 1937 2476 1943
rect 2685 1937 2716 1943
rect 2964 1937 2988 1943
rect 3101 1943 3107 1963
rect 3101 1937 3148 1943
rect 3156 1937 3164 1943
rect 3901 1937 3932 1943
rect 4324 1937 4403 1943
rect 2796 1932 2804 1936
rect 253 1917 275 1923
rect 429 1897 451 1903
rect 445 1884 451 1897
rect 493 1903 499 1923
rect 573 1917 588 1923
rect 621 1917 636 1923
rect 1853 1917 1868 1923
rect 1924 1916 1932 1924
rect 2468 1917 2483 1923
rect 2781 1917 2803 1923
rect 2861 1917 2892 1923
rect 3357 1917 3411 1923
rect 3581 1917 3603 1923
rect 3684 1916 3692 1924
rect 3748 1916 3756 1924
rect 3773 1917 3811 1923
rect 4253 1917 4284 1923
rect 484 1897 499 1903
rect 948 1897 979 1903
rect 1012 1897 1043 1903
rect 1645 1903 1651 1916
rect 1581 1897 1651 1903
rect 1933 1897 1964 1903
rect 1972 1897 1987 1903
rect 1997 1897 2012 1903
rect 3172 1897 3187 1903
rect 3444 1897 3491 1903
rect 3652 1897 3683 1903
rect 3732 1897 3747 1903
rect 4173 1897 4204 1903
rect 4669 1897 4740 1903
rect 125 1877 172 1883
rect 532 1877 547 1883
rect 580 1877 595 1883
rect 692 1877 707 1883
rect 845 1877 860 1883
rect 1524 1877 1539 1883
rect 1709 1877 1724 1883
rect 1853 1877 1891 1883
rect 1652 1856 1660 1864
rect 1853 1857 1859 1877
rect 1956 1877 1971 1883
rect 2680 1876 2684 1884
rect 2829 1877 2844 1883
rect 2877 1877 2892 1883
rect 3460 1877 3475 1883
rect 4061 1883 4067 1896
rect 4732 1892 4740 1897
rect 4909 1897 4924 1903
rect 5133 1897 5148 1903
rect 4045 1877 4067 1883
rect 4132 1877 4147 1883
rect 4973 1877 4995 1883
rect 5005 1877 5036 1883
rect 4989 1864 4995 1877
rect 5133 1877 5139 1897
rect 5357 1903 5363 1923
rect 5501 1917 5523 1923
rect 5572 1916 5580 1924
rect 5357 1897 5372 1903
rect 5581 1897 5628 1903
rect 6045 1897 6083 1903
rect 5284 1877 5315 1883
rect 5604 1877 5619 1883
rect 5692 1877 5708 1883
rect 5692 1876 5700 1877
rect 5852 1877 5868 1883
rect 5852 1876 5860 1877
rect 6008 1877 6028 1883
rect 6221 1877 6236 1883
rect 4004 1857 4028 1863
rect 4100 1856 4108 1864
rect 4317 1857 4332 1863
rect 4548 1857 4572 1863
rect 4813 1857 4828 1863
rect 5172 1856 5180 1864
rect 5412 1856 5420 1864
rect 6125 1857 6147 1863
rect 122 1836 124 1844
rect 292 1837 307 1843
rect 346 1836 348 1844
rect 506 1836 508 1844
rect 788 1836 790 1844
rect 1540 1836 1542 1844
rect 2810 1836 2812 1844
rect 3325 1837 3340 1843
rect 4445 1837 4460 1843
rect 4628 1836 4630 1844
rect 5076 1836 5080 1844
rect 3112 1806 3118 1814
rect 3126 1806 3132 1814
rect 3140 1806 3146 1814
rect 3154 1806 3160 1814
rect 2349 1777 2364 1783
rect 2440 1776 2444 1784
rect 2564 1776 2568 1784
rect 5208 1776 5212 1784
rect 5274 1776 5276 1784
rect 5762 1777 5788 1783
rect 6221 1777 6252 1783
rect 580 1757 611 1763
rect 3220 1757 3244 1763
rect 3517 1757 3555 1763
rect 3965 1757 4003 1763
rect 644 1737 659 1743
rect 781 1737 796 1743
rect 925 1737 940 1743
rect 948 1737 979 1743
rect 1741 1737 1772 1743
rect 2260 1737 2275 1743
rect 2756 1737 2771 1743
rect 2781 1737 2812 1743
rect 2852 1737 2883 1743
rect 2916 1737 2931 1743
rect 3364 1737 3411 1743
rect 420 1717 435 1723
rect 541 1717 556 1723
rect 621 1717 643 1723
rect 1117 1717 1123 1736
rect 1149 1717 1155 1736
rect 1229 1717 1244 1723
rect 1428 1717 1459 1723
rect 1476 1717 1507 1723
rect 1540 1717 1619 1723
rect 1821 1717 1859 1723
rect 317 1697 332 1703
rect 781 1697 819 1703
rect 1533 1697 1548 1703
rect 1821 1697 1827 1717
rect 2244 1717 2291 1723
rect 2653 1717 2668 1723
rect 2980 1717 2995 1723
rect 3108 1717 3171 1723
rect 3213 1717 3228 1723
rect 3348 1717 3427 1723
rect 3533 1717 3548 1723
rect 3757 1723 3763 1743
rect 3917 1737 3955 1743
rect 4372 1737 4387 1743
rect 4493 1743 4499 1763
rect 4509 1757 4547 1763
rect 4829 1744 4835 1763
rect 4484 1737 4499 1743
rect 4792 1736 4796 1744
rect 4941 1743 4947 1763
rect 4836 1737 4851 1743
rect 4909 1737 4947 1743
rect 5245 1737 5260 1743
rect 5316 1737 5331 1743
rect 3748 1717 3763 1723
rect 3789 1717 3827 1723
rect 1860 1696 1868 1704
rect 221 1677 252 1683
rect 836 1677 851 1683
rect 1949 1683 1955 1703
rect 1949 1677 1971 1683
rect 2292 1676 2294 1684
rect 2397 1683 2403 1703
rect 3293 1697 3315 1703
rect 3821 1697 3827 1717
rect 4148 1717 4179 1723
rect 4253 1717 4291 1723
rect 4253 1697 4259 1717
rect 4397 1717 4435 1723
rect 4461 1717 4476 1723
rect 4429 1697 4435 1717
rect 4596 1717 4627 1723
rect 4637 1717 4700 1723
rect 4740 1717 4756 1723
rect 4748 1712 4756 1717
rect 5021 1717 5107 1723
rect 4653 1697 4723 1703
rect 5021 1697 5027 1717
rect 5613 1717 5644 1723
rect 5661 1717 5708 1723
rect 5821 1723 5827 1743
rect 5821 1717 5852 1723
rect 5581 1697 5596 1703
rect 5874 1696 5884 1704
rect 6221 1697 6236 1703
rect 2372 1677 2403 1683
rect 2468 1677 2499 1683
rect 3060 1677 3091 1683
rect 1620 1656 1622 1664
rect 1290 1636 1292 1644
rect 1402 1636 1404 1644
rect 1508 1636 1510 1644
rect 1796 1636 1798 1644
rect 2042 1636 2044 1644
rect 3674 1636 3676 1644
rect 3850 1636 3852 1644
rect 4122 1636 4124 1644
rect 4458 1636 4460 1644
rect 4996 1636 4998 1644
rect 1560 1606 1566 1614
rect 1574 1606 1580 1614
rect 1588 1606 1594 1614
rect 1602 1606 1608 1614
rect 4632 1606 4638 1614
rect 4646 1606 4652 1614
rect 4660 1606 4666 1614
rect 4674 1606 4680 1614
rect 3194 1576 3196 1584
rect 5466 1576 5468 1584
rect 1108 1536 1110 1544
rect 1496 1536 1500 1544
rect 2797 1537 2828 1543
rect 3085 1543 3091 1563
rect 3864 1556 3868 1564
rect 3085 1537 3155 1543
rect 3149 1524 3155 1537
rect 4468 1536 4470 1544
rect 5108 1536 5110 1544
rect 5677 1537 5708 1543
rect 29 1517 67 1523
rect 164 1497 179 1503
rect 516 1497 531 1503
rect 973 1497 988 1503
rect 1092 1497 1107 1503
rect 1213 1503 1219 1523
rect 1181 1497 1219 1503
rect 1325 1503 1331 1523
rect 1757 1517 1772 1523
rect 1821 1517 1836 1523
rect 2653 1517 2675 1523
rect 3156 1517 3171 1523
rect 3533 1517 3548 1523
rect 4180 1517 4195 1523
rect 1325 1497 1340 1503
rect 1933 1503 1939 1516
rect 1885 1497 1907 1503
rect 1933 1497 1955 1503
rect 109 1477 124 1483
rect 1901 1484 1907 1497
rect 2237 1497 2275 1503
rect 2925 1497 2956 1503
rect 3492 1497 3507 1503
rect 4237 1497 4252 1503
rect 1389 1477 1404 1483
rect 125 1457 131 1476
rect 804 1457 828 1463
rect 1389 1457 1395 1477
rect 1565 1477 1596 1483
rect 1757 1477 1779 1483
rect 2148 1477 2179 1483
rect 2573 1477 2588 1483
rect 2989 1477 3004 1483
rect 3325 1477 3340 1483
rect 3453 1477 3491 1483
rect 3725 1477 3747 1483
rect 4237 1477 4243 1497
rect 4429 1497 4467 1503
rect 4596 1497 4611 1503
rect 5037 1497 5052 1503
rect 6125 1497 6140 1503
rect 4292 1477 4307 1483
rect 5373 1477 5404 1483
rect 5757 1477 5788 1483
rect 1924 1457 1948 1463
rect 2221 1457 2236 1463
rect 3677 1457 3715 1463
rect 4676 1457 4732 1463
rect 5396 1457 5411 1463
rect 5597 1457 5635 1463
rect 372 1436 374 1444
rect 442 1436 444 1444
rect 602 1436 604 1444
rect 1050 1436 1052 1444
rect 2122 1436 2124 1444
rect 2532 1436 2534 1444
rect 2621 1437 2636 1443
rect 2970 1436 2972 1444
rect 3252 1436 3254 1444
rect 3562 1436 3564 1444
rect 5218 1437 5244 1443
rect 5293 1437 5308 1443
rect 5802 1436 5804 1444
rect 6008 1436 6012 1444
rect 3112 1406 3118 1414
rect 3126 1406 3132 1414
rect 3140 1406 3146 1414
rect 3154 1406 3160 1414
rect 3300 1376 3302 1384
rect 3812 1376 3814 1384
rect 3853 1377 3868 1383
rect 5565 1377 5580 1383
rect 909 1357 924 1363
rect 4093 1357 4108 1363
rect 4244 1356 4252 1364
rect 4372 1357 4387 1363
rect 4957 1357 4979 1363
rect 5428 1357 5443 1363
rect 29 1337 67 1343
rect 541 1337 556 1343
rect 733 1337 748 1343
rect 964 1337 979 1343
rect 1044 1337 1075 1343
rect 1437 1337 1452 1343
rect 1700 1337 1715 1343
rect 1780 1337 1795 1343
rect 1869 1337 1884 1343
rect 1956 1337 1971 1343
rect 2109 1343 2115 1356
rect 2109 1337 2131 1343
rect 2173 1337 2188 1343
rect 2365 1337 2387 1343
rect 2708 1337 2739 1343
rect 2916 1337 2931 1343
rect 3101 1337 3171 1343
rect 3437 1337 3452 1343
rect 3933 1337 3964 1343
rect 4612 1337 4627 1343
rect 4644 1337 4707 1343
rect 4861 1337 4876 1343
rect 5229 1337 5260 1343
rect 5300 1337 5315 1343
rect 5437 1337 5468 1343
rect 5476 1337 5491 1343
rect 5645 1337 5692 1343
rect 5764 1337 5811 1343
rect 532 1317 579 1323
rect 797 1317 812 1323
rect 980 1317 995 1323
rect 1300 1317 1315 1323
rect 1421 1317 1468 1323
rect 605 1297 643 1303
rect 1309 1297 1315 1317
rect 1757 1317 1788 1323
rect 2068 1317 2083 1323
rect 3028 1317 3043 1323
rect 2452 1297 2467 1303
rect 3037 1297 3043 1317
rect 3981 1317 4003 1323
rect 4061 1317 4099 1323
rect 4164 1317 4179 1323
rect 4509 1317 4540 1323
rect 4573 1317 4611 1323
rect 3373 1297 3395 1303
rect 3549 1297 3571 1303
rect 3036 1284 3044 1288
rect 93 1277 108 1283
rect 189 1277 268 1283
rect 2060 1277 2083 1283
rect 3652 1276 3654 1284
rect 4429 1283 4435 1303
rect 4477 1297 4492 1303
rect 4605 1297 4611 1317
rect 4781 1317 4796 1323
rect 5421 1317 5436 1323
rect 5444 1317 5507 1323
rect 5741 1317 5772 1323
rect 5780 1317 5827 1323
rect 5837 1317 5868 1323
rect 4749 1297 4764 1303
rect 5981 1297 6012 1303
rect 4413 1277 4435 1283
rect 5508 1276 5510 1284
rect 2036 1256 2038 1264
rect 580 1236 582 1244
rect 938 1236 940 1244
rect 996 1236 998 1244
rect 1418 1236 1420 1244
rect 1476 1236 1478 1244
rect 2346 1236 2348 1244
rect 3594 1236 3596 1244
rect 3754 1236 3756 1244
rect 4346 1236 4348 1244
rect 5060 1236 5062 1244
rect 5178 1236 5180 1244
rect 1560 1206 1566 1214
rect 1574 1206 1580 1214
rect 1588 1206 1594 1214
rect 1602 1206 1608 1214
rect 4632 1206 4638 1214
rect 4646 1206 4652 1214
rect 4660 1206 4666 1214
rect 4674 1206 4680 1214
rect 1748 1176 1750 1184
rect 3117 1177 3164 1183
rect 3764 1176 3766 1184
rect 1828 1137 1891 1143
rect 2013 1143 2019 1163
rect 2013 1137 2028 1143
rect 2205 1143 2211 1163
rect 2205 1137 2220 1143
rect 2244 1137 2275 1143
rect 2349 1137 2403 1143
rect 2349 1124 2355 1137
rect 2452 1137 2467 1143
rect 2660 1137 2691 1143
rect 2932 1136 2934 1144
rect 3293 1137 3324 1143
rect 4376 1136 4380 1144
rect 5460 1136 5462 1144
rect 2684 1124 2692 1128
rect 1533 1117 1564 1123
rect 1828 1117 1843 1123
rect 2020 1117 2035 1123
rect 3021 1117 3059 1123
rect 3469 1117 3484 1123
rect 3789 1117 3811 1123
rect 5549 1117 5571 1123
rect 77 1097 108 1103
rect 333 1097 348 1103
rect 868 1097 883 1103
rect 980 1097 1011 1103
rect 1229 1097 1260 1103
rect 1316 1097 1331 1103
rect 1693 1097 1724 1103
rect 2477 1097 2499 1103
rect 2781 1097 2844 1103
rect 2852 1097 2867 1103
rect 2916 1097 2931 1103
rect 3005 1097 3036 1103
rect 3965 1097 3996 1103
rect 4141 1097 4156 1103
rect 4260 1097 4275 1103
rect 4552 1096 4556 1104
rect 116 1077 147 1083
rect 253 1077 268 1083
rect 276 1077 291 1083
rect 461 1083 467 1096
rect 461 1077 483 1083
rect 1149 1077 1164 1083
rect 1389 1077 1404 1083
rect 1629 1077 1660 1083
rect 2804 1077 2851 1083
rect 3196 1077 3212 1083
rect 3196 1076 3204 1077
rect 3828 1077 3859 1083
rect 4301 1077 4323 1083
rect 4301 1064 4307 1077
rect 4701 1083 4707 1103
rect 5213 1097 5228 1103
rect 5421 1097 5459 1103
rect 5693 1097 5708 1103
rect 5796 1096 5800 1104
rect 4596 1077 4611 1083
rect 4621 1077 4707 1083
rect 2788 1057 2803 1063
rect 3380 1056 3388 1064
rect 3636 1056 3644 1064
rect 3885 1057 3900 1063
rect 4244 1057 4268 1063
rect 4605 1057 4611 1077
rect 4765 1077 4803 1083
rect 5165 1077 5187 1083
rect 5384 1077 5404 1083
rect 5741 1083 5747 1096
rect 5741 1077 5763 1083
rect 292 1036 294 1044
rect 612 1036 614 1044
rect 778 1036 780 1044
rect 1501 1037 1516 1043
rect 3140 1037 3164 1043
rect 3508 1036 3510 1044
rect 5064 1036 5068 1044
rect 5588 1037 5603 1043
rect 3112 1006 3118 1014
rect 3126 1006 3132 1014
rect 3140 1006 3146 1014
rect 3154 1006 3160 1014
rect 1869 977 1884 983
rect 1933 977 1948 983
rect 2984 976 2988 984
rect 3053 977 3100 983
rect 4296 976 4300 984
rect 4362 976 4364 984
rect 5284 976 5288 984
rect 2068 956 2076 964
rect 173 937 188 943
rect 340 937 355 943
rect 1204 937 1235 943
rect 1709 937 1724 943
rect 1832 936 1836 944
rect 2269 937 2284 943
rect 2868 937 2883 943
rect 2893 937 2931 943
rect 3213 937 3228 943
rect 3501 937 3516 943
rect 3533 937 3564 943
rect 3645 943 3651 963
rect 3716 957 3731 963
rect 4077 957 4115 963
rect 4413 957 4435 963
rect 4445 957 4460 963
rect 4829 957 4860 963
rect 3645 937 3676 943
rect 4109 937 4147 943
rect 4413 937 4428 943
rect 4493 937 4524 943
rect 4564 937 4588 943
rect 4813 937 4844 943
rect 4932 937 4947 943
rect 5421 943 5427 963
rect 5412 937 5427 943
rect 5501 943 5507 963
rect 5501 937 5516 943
rect 5725 943 5731 963
rect 5693 937 5731 943
rect 1213 917 1228 923
rect 1245 917 1283 923
rect 509 897 524 903
rect 628 897 659 903
rect 948 897 963 903
rect 1053 897 1068 903
rect 1277 897 1283 917
rect 1549 917 1612 923
rect 1645 917 1683 923
rect 1485 897 1523 903
rect 1540 896 1548 904
rect 1677 897 1683 917
rect 2253 917 2300 923
rect 2516 917 2532 923
rect 2524 912 2532 917
rect 3220 917 3251 923
rect 3284 917 3315 923
rect 3412 917 3427 923
rect 3501 917 3523 923
rect 3501 904 3507 917
rect 3597 917 3612 923
rect 4637 917 4684 923
rect 4740 917 4771 923
rect 5757 917 5779 923
rect 6100 917 6115 923
rect 1892 897 1907 903
rect 2077 897 2092 903
rect 2525 897 2540 903
rect 292 877 307 883
rect 877 877 931 883
rect 1028 877 1043 883
rect 1380 877 1436 883
rect 1933 877 1948 883
rect 2365 877 2396 883
rect 2660 876 2662 884
rect 2813 883 2819 903
rect 3277 897 3292 903
rect 3325 897 3347 903
rect 3613 897 3635 903
rect 4189 897 4211 903
rect 2813 877 2835 883
rect 3901 877 3916 883
rect 5386 876 5388 884
rect 826 836 828 844
rect 2250 836 2252 844
rect 2842 836 2844 844
rect 3176 836 3180 844
rect 6036 836 6040 844
rect 1560 806 1566 814
rect 1574 806 1580 814
rect 1588 806 1594 814
rect 1602 806 1608 814
rect 4632 806 4638 814
rect 4646 806 4652 814
rect 4660 806 4666 814
rect 4674 806 4680 814
rect 660 776 662 784
rect 2186 776 2188 784
rect 5050 776 5052 784
rect 6212 776 6214 784
rect 420 736 422 744
rect 2148 736 2150 744
rect 4980 736 4982 744
rect 980 717 995 723
rect 1076 716 1084 724
rect 1924 717 1939 723
rect 2045 717 2060 723
rect 3117 717 3187 723
rect 3389 717 3404 723
rect 4429 717 4444 723
rect 180 697 227 703
rect 404 697 419 703
rect 685 703 691 716
rect 685 697 707 703
rect 877 697 892 703
rect 973 697 988 703
rect 189 677 204 683
rect 557 677 588 683
rect 749 677 780 683
rect 973 677 979 697
rect 1021 697 1068 703
rect 1661 697 1731 703
rect 2301 697 2332 703
rect 2660 697 2739 703
rect 3005 697 3020 703
rect 3076 697 3091 703
rect 3101 697 3164 703
rect 3629 697 3660 703
rect 3740 703 3748 708
rect 3740 697 3763 703
rect 3837 697 3875 703
rect 3885 697 3916 703
rect 4349 697 4364 703
rect 4484 697 4499 703
rect 4717 697 4732 703
rect 4812 703 4820 708
rect 4812 697 4828 703
rect 4941 697 4979 703
rect 5277 697 5292 703
rect 5356 703 5364 708
rect 5356 697 5372 703
rect 5421 697 5459 703
rect 5828 696 5832 704
rect 5892 697 5907 703
rect 6013 697 6028 703
rect 1044 677 1059 683
rect 1172 677 1203 683
rect 1357 677 1388 683
rect 1460 677 1491 683
rect 2253 677 2268 683
rect 84 657 99 663
rect 596 656 604 664
rect 788 656 796 664
rect 1421 657 1443 663
rect 1576 657 1651 663
rect 2253 657 2259 677
rect 2349 677 2364 683
rect 2676 677 2723 683
rect 3037 677 3068 683
rect 3204 677 3235 683
rect 3245 677 3260 683
rect 3396 677 3411 683
rect 3421 677 3452 683
rect 3604 677 3619 683
rect 4221 677 4243 683
rect 4500 677 4515 683
rect 4780 677 4796 683
rect 4780 676 4788 677
rect 4845 677 4867 683
rect 5389 677 5411 683
rect 5421 677 5452 683
rect 2573 657 2604 663
rect 2685 657 2700 663
rect 2824 656 2828 664
rect 3597 657 3603 676
rect 132 637 147 643
rect 906 636 908 644
rect 954 636 956 644
rect 1746 637 1772 643
rect 2404 636 2406 644
rect 3300 637 3315 643
rect 4088 636 4092 644
rect 5108 636 5110 644
rect 5498 636 5500 644
rect 5576 636 5580 644
rect 3112 606 3118 614
rect 3126 606 3132 614
rect 3140 606 3146 614
rect 3154 606 3160 614
rect 1341 577 1356 583
rect 1549 577 1596 583
rect 1661 577 1676 583
rect 1725 577 1740 583
rect 2260 576 2262 584
rect 2344 576 2348 584
rect 2420 576 2422 584
rect 2680 576 2684 584
rect 2756 576 2758 584
rect 3444 576 3446 584
rect 3576 576 3580 584
rect 4776 576 4780 584
rect 1181 557 1203 563
rect 2829 557 2844 563
rect 3725 557 3747 563
rect 173 537 188 543
rect 388 537 403 543
rect 772 537 787 543
rect 77 517 147 523
rect 189 517 212 523
rect 204 512 212 517
rect 372 517 419 523
rect 756 517 803 523
rect 909 523 915 543
rect 1304 536 1308 544
rect 1492 537 1523 543
rect 2061 543 2067 556
rect 2061 537 2083 543
rect 2077 524 2083 537
rect 2589 537 2604 543
rect 2868 537 2883 543
rect 3053 537 3116 543
rect 3229 537 3244 543
rect 3709 537 3724 543
rect 3741 543 3747 557
rect 4964 557 4979 563
rect 4989 557 5011 563
rect 3741 537 3763 543
rect 3869 537 3884 543
rect 3917 537 3932 543
rect 4164 537 4179 543
rect 4644 537 4707 543
rect 4829 537 4844 543
rect 5005 543 5011 557
rect 5421 557 5443 563
rect 5869 557 5884 563
rect 5005 537 5027 543
rect 5709 537 5731 543
rect 884 517 915 523
rect 2205 517 2220 523
rect 2829 517 2876 523
rect 1092 497 1107 503
rect 1149 497 1164 503
rect 420 476 422 484
rect 1389 483 1395 503
rect 2477 497 2499 503
rect 2829 497 2835 517
rect 2948 517 2979 523
rect 3453 517 3491 523
rect 3362 496 3372 504
rect 3453 497 3459 517
rect 3700 517 3779 523
rect 3805 517 3836 523
rect 3805 497 3811 517
rect 3876 517 3891 523
rect 4093 517 4124 523
rect 4525 517 4579 523
rect 4964 517 5043 523
rect 5229 517 5267 523
rect 5373 517 5388 523
rect 5677 517 5692 523
rect 5885 517 5907 523
rect 5997 517 6028 523
rect 4125 497 4131 516
rect 4573 497 4611 503
rect 4724 497 4739 503
rect 5293 497 5331 503
rect 5389 497 5404 503
rect 1364 477 1395 483
rect 3156 477 3180 483
rect 4196 476 4198 484
rect 5549 477 5580 483
rect 932 436 934 444
rect 5268 436 5270 444
rect 1560 406 1566 414
rect 1574 406 1580 414
rect 1588 406 1594 414
rect 1602 406 1608 414
rect 4632 406 4638 414
rect 4646 406 4652 414
rect 4660 406 4666 414
rect 4674 406 4680 414
rect 804 376 806 384
rect 1930 376 1932 384
rect 2024 376 2028 384
rect 2890 376 2892 384
rect 2964 376 2968 384
rect 3690 376 3692 384
rect 4548 376 4550 384
rect 5108 376 5110 384
rect 5866 376 5868 384
rect 6052 376 6056 384
rect 29 337 60 343
rect 1405 337 1436 343
rect 1405 317 1411 337
rect 1834 336 1836 344
rect 2712 336 2716 344
rect 3428 336 3432 344
rect 5412 337 5443 343
rect 5924 337 5939 343
rect 1796 317 1811 323
rect 893 297 908 303
rect 916 297 931 303
rect 941 297 972 303
rect 1757 297 1779 303
rect 2221 297 2236 303
rect 2413 303 2419 323
rect 4381 317 4403 323
rect 5172 316 5180 324
rect 5828 317 5843 323
rect 2269 297 2307 303
rect 2317 297 2387 303
rect 2413 297 2460 303
rect 2621 297 2652 303
rect 3069 297 3107 303
rect 3549 297 3571 303
rect 3604 297 3619 303
rect 3629 297 3660 303
rect 4077 297 4092 303
rect 4148 297 4163 303
rect 4205 297 4268 303
rect 685 277 700 283
rect 349 257 364 263
rect 685 257 691 277
rect 1272 276 1276 284
rect 1368 276 1372 284
rect 1956 277 1971 283
rect 2173 277 2188 283
rect 2413 277 2428 283
rect 2468 277 2499 283
rect 2525 277 2547 283
rect 3021 277 3059 283
rect 3156 277 3171 283
rect 3213 277 3228 283
rect 3716 277 3731 283
rect 4036 277 4051 283
rect 4157 277 4163 297
rect 4509 297 4547 303
rect 4788 297 4803 303
rect 5181 297 5196 303
rect 5204 297 5267 303
rect 5288 297 5324 303
rect 4276 277 4291 283
rect 4413 277 4428 283
rect 724 257 748 263
rect 2205 257 2243 263
rect 3076 257 3091 263
rect 3597 257 3635 263
rect 3828 257 3859 263
rect 4029 257 4051 263
rect 4413 257 4419 277
rect 5197 277 5244 283
rect 5716 257 5731 263
rect 5988 256 5996 264
rect 228 237 243 243
rect 3288 236 3292 244
rect 4644 237 4691 243
rect 5560 236 5564 244
rect 3112 206 3118 214
rect 3126 206 3132 214
rect 3140 206 3146 214
rect 3154 206 3160 214
rect 845 177 860 183
rect 1800 176 1804 184
rect 2296 176 2300 184
rect 3524 176 3526 184
rect 3608 176 3612 184
rect 3674 176 3676 184
rect 4008 176 4012 184
rect 4152 176 4156 184
rect 5421 177 5436 183
rect 5546 176 5548 184
rect 5956 176 5958 184
rect 109 143 115 163
rect 1069 157 1091 163
rect 1421 157 1436 163
rect 1956 156 1964 164
rect 2701 157 2716 163
rect 2852 157 2867 163
rect 93 123 99 143
rect 109 137 140 143
rect 93 117 108 123
rect 116 117 163 123
rect 269 123 275 143
rect 461 143 467 156
rect 429 137 467 143
rect 477 137 508 143
rect 973 137 988 143
rect 1028 137 1043 143
rect 1172 137 1187 143
rect 1229 137 1260 143
rect 1348 137 1363 143
rect 1444 137 1459 143
rect 1517 137 1532 143
rect 1837 137 1859 143
rect 1901 137 1916 143
rect 2013 137 2044 143
rect 2061 137 2099 143
rect 2196 137 2211 143
rect 2397 137 2435 143
rect 244 117 275 123
rect 1005 117 1027 123
rect 1156 117 1203 123
rect 1341 117 1356 123
rect 1437 117 1452 123
rect 1741 123 1747 136
rect 2541 137 2563 143
rect 2596 137 2627 143
rect 2660 137 2691 143
rect 2708 137 2739 143
rect 3005 143 3011 163
rect 2820 137 2835 143
rect 3005 137 3020 143
rect 3060 137 3075 143
rect 3213 143 3219 163
rect 3252 157 3283 163
rect 3133 137 3203 143
rect 3213 137 3228 143
rect 1533 117 1555 123
rect 1688 117 1747 123
rect 2157 117 2188 123
rect 2628 117 2643 123
rect 3133 123 3139 137
rect 3325 137 3363 143
rect 3460 137 3475 143
rect 3741 143 3747 163
rect 3780 156 3788 164
rect 4436 156 4444 164
rect 5156 157 5171 163
rect 5181 157 5196 163
rect 5236 157 5251 163
rect 5652 157 5667 163
rect 3741 137 3756 143
rect 3796 137 3811 143
rect 3917 137 3955 143
rect 4052 137 4067 143
rect 4189 137 4243 143
rect 4372 137 4403 143
rect 5037 137 5052 143
rect 5092 137 5123 143
rect 5508 137 5523 143
rect 5789 137 5827 143
rect 6180 137 6195 143
rect 3101 117 3139 123
rect 3220 117 3251 123
rect 3293 117 3308 123
rect 3421 117 3452 123
rect 3725 117 3740 123
rect 3773 117 3811 123
rect 52 98 56 106
rect 893 83 899 103
rect 3805 97 3811 117
rect 3885 117 3907 123
rect 4333 117 4355 123
rect 4413 117 4435 123
rect 4429 97 4435 117
rect 4877 117 4892 123
rect 4909 117 4947 123
rect 4941 97 4947 117
rect 5085 117 5107 123
rect 5085 104 5091 117
rect 5325 117 5340 123
rect 5373 117 5388 123
rect 5476 117 5507 123
rect 5668 117 5699 123
rect 5880 117 5932 123
rect 4957 97 4972 103
rect 5293 97 5308 103
rect 4428 84 4436 88
rect 852 77 899 83
rect 5370 76 5372 84
rect 292 56 294 64
rect 1560 6 1566 14
rect 1574 6 1580 14
rect 1588 6 1594 14
rect 1602 6 1608 14
rect 4632 6 4638 14
rect 4646 6 4652 14
rect 4660 6 4666 14
rect 4674 6 4680 14
<< m2contact >>
rect 3118 5806 3126 5814
rect 3132 5806 3140 5814
rect 3146 5806 3154 5814
rect 1292 5776 1300 5784
rect 1836 5776 1844 5784
rect 4908 5776 4916 5784
rect 5628 5776 5636 5784
rect 6140 5776 6148 5784
rect 124 5756 132 5764
rect 156 5756 164 5764
rect 284 5756 292 5764
rect 492 5756 500 5764
rect 508 5756 516 5764
rect 908 5756 916 5764
rect 924 5756 932 5764
rect 956 5756 964 5764
rect 1148 5756 1156 5764
rect 1212 5756 1220 5764
rect 1388 5756 1396 5764
rect 1500 5756 1508 5764
rect 1596 5756 1604 5764
rect 1676 5756 1684 5764
rect 1852 5756 1860 5764
rect 1932 5756 1940 5764
rect 1996 5756 2004 5764
rect 2348 5756 2356 5764
rect 2652 5756 2660 5764
rect 2668 5756 2676 5764
rect 2780 5756 2788 5764
rect 92 5736 100 5744
rect 124 5736 132 5744
rect 252 5736 260 5744
rect 300 5736 308 5744
rect 364 5736 372 5744
rect 396 5736 404 5744
rect 540 5736 548 5744
rect 588 5736 596 5744
rect 652 5736 660 5744
rect 668 5736 676 5744
rect 44 5716 52 5724
rect 76 5716 84 5724
rect 204 5716 212 5724
rect 236 5716 244 5724
rect 444 5716 452 5724
rect 540 5716 548 5724
rect 572 5716 580 5724
rect 588 5716 596 5724
rect 780 5736 788 5744
rect 988 5736 996 5744
rect 844 5716 852 5724
rect 1068 5736 1076 5744
rect 1116 5736 1124 5744
rect 1196 5736 1204 5744
rect 1324 5736 1332 5744
rect 1340 5736 1348 5744
rect 1468 5736 1476 5744
rect 1516 5736 1524 5744
rect 1820 5736 1828 5744
rect 1868 5736 1876 5744
rect 1932 5736 1940 5744
rect 1964 5736 1972 5744
rect 2076 5736 2084 5744
rect 2124 5736 2132 5744
rect 2140 5736 2148 5744
rect 2204 5736 2212 5744
rect 2428 5736 2436 5744
rect 2540 5736 2548 5744
rect 2700 5736 2708 5744
rect 2716 5736 2724 5744
rect 2796 5736 2804 5744
rect 2924 5736 2932 5744
rect 3020 5736 3028 5744
rect 3132 5736 3140 5744
rect 3260 5736 3268 5744
rect 3292 5736 3300 5744
rect 3548 5756 3556 5764
rect 3628 5756 3636 5764
rect 3692 5756 3700 5764
rect 3836 5756 3844 5764
rect 3932 5756 3940 5764
rect 4060 5756 4068 5764
rect 4124 5756 4132 5764
rect 4140 5756 4148 5764
rect 4172 5756 4180 5764
rect 4364 5756 4372 5764
rect 4444 5756 4452 5764
rect 4572 5756 4580 5764
rect 4588 5756 4596 5764
rect 4748 5756 4756 5764
rect 1020 5716 1028 5724
rect 1052 5716 1060 5724
rect 1388 5716 1396 5724
rect 1644 5716 1652 5724
rect 1772 5716 1780 5724
rect 1804 5716 1812 5724
rect 1932 5716 1940 5724
rect 1948 5716 1956 5724
rect 2028 5716 2036 5724
rect 2092 5716 2100 5724
rect 2156 5716 2164 5724
rect 2220 5716 2228 5724
rect 2284 5716 2292 5724
rect 2332 5716 2340 5724
rect 2380 5716 2388 5724
rect 2572 5716 2580 5724
rect 2620 5716 2628 5724
rect 2748 5716 2756 5724
rect 2812 5716 2820 5724
rect 2876 5716 2884 5724
rect 3084 5716 3092 5724
rect 3228 5716 3236 5724
rect 3516 5736 3524 5744
rect 3612 5736 3620 5744
rect 3804 5736 3812 5744
rect 4124 5736 4132 5744
rect 4220 5736 4228 5744
rect 4236 5736 4244 5744
rect 4444 5736 4452 5744
rect 4716 5736 4724 5744
rect 4764 5736 4772 5744
rect 4876 5756 4884 5764
rect 4892 5756 4900 5764
rect 4924 5756 4932 5764
rect 4988 5756 4996 5764
rect 5004 5756 5012 5764
rect 5228 5756 5236 5764
rect 5356 5756 5364 5764
rect 5452 5756 5460 5764
rect 5580 5756 5588 5764
rect 5596 5756 5604 5764
rect 5916 5756 5924 5764
rect 5996 5756 6004 5764
rect 4972 5736 4980 5744
rect 5148 5736 5156 5744
rect 5244 5736 5252 5744
rect 5452 5736 5460 5744
rect 5836 5736 5844 5744
rect 5900 5736 5908 5744
rect 6236 5736 6244 5744
rect 3420 5716 3428 5724
rect 3468 5716 3476 5724
rect 3516 5716 3524 5724
rect 60 5696 68 5704
rect 220 5696 228 5704
rect 348 5696 356 5704
rect 364 5696 372 5704
rect 396 5696 404 5704
rect 460 5696 468 5704
rect 540 5696 548 5704
rect 604 5696 612 5704
rect 812 5696 820 5704
rect 828 5696 836 5704
rect 956 5696 964 5704
rect 1052 5696 1060 5704
rect 1100 5696 1108 5704
rect 1148 5696 1156 5704
rect 1372 5696 1380 5704
rect 1420 5696 1428 5704
rect 1548 5696 1556 5704
rect 1724 5696 1732 5704
rect 1788 5696 1796 5704
rect 1900 5696 1908 5704
rect 2012 5696 2020 5704
rect 2124 5696 2132 5704
rect 2188 5696 2196 5704
rect 2252 5696 2260 5704
rect 2268 5696 2276 5704
rect 2364 5696 2372 5704
rect 2492 5696 2500 5704
rect 2572 5696 2580 5704
rect 2652 5696 2660 5704
rect 2684 5696 2692 5704
rect 2780 5696 2788 5704
rect 2860 5696 2868 5704
rect 2988 5696 2996 5704
rect 3244 5696 3252 5704
rect 3292 5696 3300 5704
rect 3340 5696 3348 5704
rect 3356 5696 3364 5704
rect 3404 5696 3412 5704
rect 3548 5696 3556 5704
rect 3580 5716 3588 5724
rect 3596 5716 3604 5724
rect 3884 5716 3892 5724
rect 3932 5716 3940 5724
rect 4188 5716 4196 5724
rect 4396 5716 4404 5724
rect 4508 5716 4516 5724
rect 4604 5716 4612 5724
rect 4684 5716 4692 5724
rect 4732 5716 4740 5724
rect 4956 5716 4964 5724
rect 5036 5716 5044 5724
rect 5068 5716 5076 5724
rect 5116 5716 5124 5724
rect 5164 5716 5172 5724
rect 5404 5716 5412 5724
rect 5516 5716 5524 5724
rect 5612 5716 5620 5724
rect 5660 5716 5668 5724
rect 5804 5718 5812 5726
rect 5916 5716 5924 5724
rect 5996 5718 6004 5726
rect 6044 5716 6052 5724
rect 6172 5716 6180 5724
rect 6220 5716 6228 5724
rect 3852 5696 3860 5704
rect 4428 5696 4436 5704
rect 4524 5696 4532 5704
rect 4844 5696 4852 5704
rect 5020 5696 5028 5704
rect 5132 5696 5140 5704
rect 5436 5696 5444 5704
rect 5532 5696 5540 5704
rect 5868 5696 5876 5704
rect 6188 5696 6196 5704
rect 28 5676 36 5684
rect 188 5676 196 5684
rect 860 5676 868 5684
rect 892 5676 900 5684
rect 972 5676 980 5684
rect 1708 5676 1716 5684
rect 1756 5676 1764 5684
rect 1884 5676 1892 5684
rect 2028 5676 2036 5684
rect 2044 5676 2052 5684
rect 2060 5676 2068 5684
rect 2300 5676 2308 5684
rect 2396 5676 2404 5684
rect 2604 5676 2612 5684
rect 3212 5676 3220 5684
rect 3388 5676 3396 5684
rect 4812 5676 4820 5684
rect 5052 5676 5060 5684
rect 5100 5676 5108 5684
rect 5676 5676 5684 5684
rect 6124 5676 6132 5684
rect 316 5656 324 5664
rect 844 5656 852 5664
rect 1772 5656 1780 5664
rect 44 5636 52 5644
rect 204 5636 212 5644
rect 732 5636 740 5644
rect 940 5636 948 5644
rect 1020 5636 1028 5644
rect 1164 5636 1172 5644
rect 1404 5636 1412 5644
rect 1452 5636 1460 5644
rect 2156 5636 2164 5644
rect 2220 5636 2228 5644
rect 2284 5636 2292 5644
rect 2380 5636 2388 5644
rect 2620 5636 2628 5644
rect 2700 5636 2708 5644
rect 2908 5636 2916 5644
rect 3228 5636 3236 5644
rect 3276 5636 3284 5644
rect 3324 5636 3332 5644
rect 3452 5636 3460 5644
rect 3740 5636 3748 5644
rect 3884 5636 3892 5644
rect 4284 5636 4292 5644
rect 4396 5636 4404 5644
rect 4860 5636 4868 5644
rect 5084 5636 5092 5644
rect 5164 5636 5172 5644
rect 5276 5636 5284 5644
rect 5404 5636 5412 5644
rect 5932 5636 5940 5644
rect 6220 5636 6228 5644
rect 1566 5606 1574 5614
rect 1580 5606 1588 5614
rect 1594 5606 1602 5614
rect 4638 5606 4646 5614
rect 4652 5606 4660 5614
rect 4666 5606 4674 5614
rect 76 5576 84 5584
rect 140 5576 148 5584
rect 284 5576 292 5584
rect 1212 5576 1220 5584
rect 1292 5576 1300 5584
rect 1548 5576 1556 5584
rect 2364 5576 2372 5584
rect 2604 5576 2612 5584
rect 4092 5576 4100 5584
rect 4268 5576 4276 5584
rect 4556 5576 4564 5584
rect 4796 5576 4804 5584
rect 5036 5576 5044 5584
rect 5356 5576 5364 5584
rect 6060 5576 6068 5584
rect 6140 5576 6148 5584
rect 780 5556 788 5564
rect 2860 5556 2868 5564
rect 3436 5556 3444 5564
rect 4908 5556 4916 5564
rect 5596 5556 5604 5564
rect 5932 5556 5940 5564
rect 92 5536 100 5544
rect 236 5536 244 5544
rect 300 5536 308 5544
rect 764 5536 772 5544
rect 1356 5536 1364 5544
rect 2156 5536 2164 5544
rect 2220 5536 2228 5544
rect 2876 5536 2884 5544
rect 2972 5536 2980 5544
rect 3260 5536 3268 5544
rect 3452 5536 3460 5544
rect 4220 5536 4228 5544
rect 4252 5536 4260 5544
rect 4604 5536 4612 5544
rect 4732 5536 4740 5544
rect 4892 5536 4900 5544
rect 5020 5536 5028 5544
rect 5292 5536 5300 5544
rect 5468 5536 5476 5544
rect 5484 5536 5492 5544
rect 5516 5536 5524 5544
rect 6076 5536 6084 5544
rect 44 5516 52 5524
rect 60 5516 68 5524
rect 204 5516 212 5524
rect 268 5516 276 5524
rect 732 5516 740 5524
rect 1052 5516 1060 5524
rect 1100 5516 1108 5524
rect 1324 5516 1332 5524
rect 1372 5516 1380 5524
rect 1436 5516 1444 5524
rect 1452 5516 1460 5524
rect 1692 5516 1700 5524
rect 1932 5516 1940 5524
rect 2108 5516 2116 5524
rect 2124 5516 2132 5524
rect 2188 5516 2196 5524
rect 2284 5516 2292 5524
rect 2428 5516 2436 5524
rect 2652 5516 2660 5524
rect 2940 5516 2948 5524
rect 2988 5516 2996 5524
rect 3116 5516 3124 5524
rect 3292 5516 3300 5524
rect 3340 5516 3348 5524
rect 3420 5516 3428 5524
rect 3628 5516 3636 5524
rect 3932 5516 3940 5524
rect 3964 5516 3972 5524
rect 4156 5516 4164 5524
rect 4284 5516 4292 5524
rect 4300 5516 4308 5524
rect 4492 5516 4500 5524
rect 4524 5516 4532 5524
rect 4636 5516 4644 5524
rect 4700 5516 4708 5524
rect 4924 5516 4932 5524
rect 5052 5516 5060 5524
rect 5340 5516 5348 5524
rect 5436 5516 5444 5524
rect 5548 5516 5556 5524
rect 5564 5516 5572 5524
rect 5676 5516 5684 5524
rect 5692 5516 5700 5524
rect 5788 5516 5796 5524
rect 5836 5516 5844 5524
rect 44 5496 52 5504
rect 76 5496 84 5504
rect 140 5496 148 5504
rect 172 5496 180 5504
rect 236 5496 244 5504
rect 284 5496 292 5504
rect 348 5496 356 5504
rect 380 5496 388 5504
rect 412 5496 420 5504
rect 428 5496 436 5504
rect 492 5496 500 5504
rect 668 5496 676 5504
rect 748 5496 756 5504
rect 876 5496 884 5504
rect 908 5496 916 5504
rect 956 5496 964 5504
rect 988 5496 996 5504
rect 1100 5496 1108 5504
rect 1292 5496 1300 5504
rect 1404 5496 1412 5504
rect 1420 5496 1428 5504
rect 1500 5496 1508 5504
rect 1612 5496 1620 5504
rect 1724 5496 1732 5504
rect 1756 5496 1764 5504
rect 1884 5496 1892 5504
rect 1916 5496 1924 5504
rect 2140 5496 2148 5504
rect 2172 5496 2180 5504
rect 2204 5496 2212 5504
rect 2396 5496 2404 5504
rect 2412 5496 2420 5504
rect 2636 5496 2644 5504
rect 2668 5496 2676 5504
rect 2748 5496 2756 5504
rect 2764 5496 2772 5504
rect 2860 5496 2868 5504
rect 2956 5496 2964 5504
rect 3004 5496 3012 5504
rect 3228 5496 3236 5504
rect 3276 5496 3284 5504
rect 3404 5496 3412 5504
rect 3436 5496 3444 5504
rect 3708 5496 3716 5504
rect 4044 5496 4052 5504
rect 4108 5496 4116 5504
rect 4268 5496 4276 5504
rect 4316 5496 4324 5504
rect 4332 5496 4340 5504
rect 4604 5496 4612 5504
rect 4716 5496 4724 5504
rect 4748 5496 4756 5504
rect 4908 5496 4916 5504
rect 4940 5496 4948 5504
rect 5036 5496 5044 5504
rect 5068 5496 5076 5504
rect 5100 5496 5108 5504
rect 5132 5496 5140 5504
rect 5212 5496 5220 5504
rect 5372 5496 5380 5504
rect 5452 5496 5460 5504
rect 5532 5496 5540 5504
rect 5596 5496 5604 5504
rect 5708 5496 5716 5504
rect 5868 5496 5876 5504
rect 5916 5496 5924 5504
rect 5996 5496 6004 5504
rect 6060 5496 6068 5504
rect 6108 5496 6116 5504
rect 6156 5496 6164 5504
rect 6236 5496 6244 5504
rect 12 5476 20 5484
rect 124 5476 132 5484
rect 188 5476 196 5484
rect 252 5476 260 5484
rect 332 5476 340 5484
rect 396 5476 404 5484
rect 444 5476 452 5484
rect 508 5476 516 5484
rect 604 5476 612 5484
rect 620 5476 628 5484
rect 716 5476 724 5484
rect 796 5476 804 5484
rect 1004 5476 1012 5484
rect 1260 5476 1268 5484
rect 1276 5476 1284 5484
rect 1340 5476 1348 5484
rect 1388 5476 1396 5484
rect 1484 5476 1492 5484
rect 1516 5476 1524 5484
rect 1660 5476 1668 5484
rect 1708 5476 1716 5484
rect 1772 5476 1780 5484
rect 1868 5476 1876 5484
rect 1980 5476 1988 5484
rect 2044 5476 2052 5484
rect 2092 5476 2100 5484
rect 2284 5476 2292 5484
rect 2332 5476 2340 5484
rect 2380 5476 2388 5484
rect 2444 5476 2452 5484
rect 2540 5476 2548 5484
rect 2572 5476 2580 5484
rect 2620 5476 2628 5484
rect 2652 5476 2660 5484
rect 2684 5476 2692 5484
rect 2716 5476 2724 5484
rect 2732 5476 2740 5484
rect 3020 5476 3028 5484
rect 3068 5476 3076 5484
rect 3180 5476 3188 5484
rect 3212 5476 3220 5484
rect 3276 5476 3284 5484
rect 3308 5476 3316 5484
rect 3388 5476 3396 5484
rect 3484 5476 3492 5484
rect 3596 5476 3604 5484
rect 3724 5476 3732 5484
rect 3772 5476 3780 5484
rect 3868 5476 3876 5484
rect 3884 5476 3892 5484
rect 3932 5476 3940 5484
rect 3980 5476 3988 5484
rect 3996 5476 4004 5484
rect 4060 5476 4068 5484
rect 4092 5476 4100 5484
rect 4124 5476 4132 5484
rect 4156 5476 4164 5484
rect 4188 5480 4196 5488
rect 4364 5476 4372 5484
rect 4492 5476 4500 5484
rect 4588 5476 4596 5484
rect 4764 5476 4772 5484
rect 4860 5476 4868 5484
rect 4956 5476 4964 5484
rect 5084 5476 5092 5484
rect 5116 5476 5124 5484
rect 5196 5476 5204 5484
rect 5228 5476 5236 5484
rect 5388 5476 5396 5484
rect 5612 5476 5620 5484
rect 5676 5476 5684 5484
rect 5788 5476 5796 5484
rect 5804 5476 5812 5484
rect 5900 5476 5908 5484
rect 6172 5476 6180 5484
rect 6252 5476 6260 5484
rect 444 5456 452 5464
rect 460 5456 468 5464
rect 796 5456 804 5464
rect 908 5456 916 5464
rect 940 5456 948 5464
rect 988 5456 996 5464
rect 1116 5456 1124 5464
rect 1148 5456 1156 5464
rect 1644 5456 1652 5464
rect 1916 5456 1924 5464
rect 1996 5456 2004 5464
rect 2092 5456 2100 5464
rect 2348 5456 2356 5464
rect 2556 5456 2564 5464
rect 2716 5456 2724 5464
rect 2812 5456 2820 5464
rect 2828 5456 2836 5464
rect 2924 5456 2932 5464
rect 3052 5456 3060 5464
rect 3180 5456 3188 5464
rect 3356 5456 3364 5464
rect 3724 5456 3732 5464
rect 3980 5456 3988 5464
rect 4156 5456 4164 5464
rect 4380 5456 4388 5464
rect 4572 5456 4580 5464
rect 4972 5456 4980 5464
rect 4988 5456 4996 5464
rect 5244 5456 5252 5464
rect 5340 5456 5348 5464
rect 5404 5456 5412 5464
rect 5420 5456 5428 5464
rect 5916 5456 5924 5464
rect 5948 5456 5956 5464
rect 6012 5456 6020 5464
rect 380 5436 388 5444
rect 540 5436 548 5444
rect 1132 5436 1140 5444
rect 1468 5436 1476 5444
rect 1676 5436 1684 5444
rect 1756 5436 1764 5444
rect 1900 5436 1908 5444
rect 2268 5436 2276 5444
rect 2316 5436 2324 5444
rect 2508 5436 2516 5444
rect 2796 5436 2804 5444
rect 2908 5436 2916 5444
rect 2972 5436 2980 5444
rect 3196 5436 3204 5444
rect 3324 5436 3332 5444
rect 3372 5436 3380 5444
rect 3532 5436 3540 5444
rect 3644 5436 3652 5444
rect 3692 5436 3700 5444
rect 3804 5436 3812 5444
rect 3916 5436 3924 5444
rect 5516 5436 5524 5444
rect 6188 5436 6196 5444
rect 3118 5406 3126 5414
rect 3132 5406 3140 5414
rect 3146 5406 3154 5414
rect 124 5376 132 5384
rect 204 5376 212 5384
rect 268 5376 276 5384
rect 348 5376 356 5384
rect 444 5376 452 5384
rect 588 5376 596 5384
rect 652 5376 660 5384
rect 764 5376 772 5384
rect 1004 5376 1012 5384
rect 1148 5376 1156 5384
rect 1948 5376 1956 5384
rect 2092 5376 2100 5384
rect 2220 5376 2228 5384
rect 2300 5376 2308 5384
rect 2428 5376 2436 5384
rect 2572 5376 2580 5384
rect 2828 5376 2836 5384
rect 3596 5376 3604 5384
rect 3948 5376 3956 5384
rect 4060 5376 4068 5384
rect 4108 5376 4116 5384
rect 4332 5376 4340 5384
rect 4428 5376 4436 5384
rect 4588 5376 4596 5384
rect 4700 5376 4708 5384
rect 4780 5376 4788 5384
rect 4956 5376 4964 5384
rect 5052 5376 5060 5384
rect 5116 5376 5124 5384
rect 5404 5376 5412 5384
rect 5612 5376 5620 5384
rect 5724 5376 5732 5384
rect 5916 5376 5924 5384
rect 5980 5376 5988 5384
rect 6172 5376 6180 5384
rect 6204 5376 6212 5384
rect 140 5356 148 5364
rect 220 5356 228 5364
rect 492 5356 500 5364
rect 604 5356 612 5364
rect 844 5356 852 5364
rect 1068 5356 1076 5364
rect 1532 5356 1540 5364
rect 1692 5356 1700 5364
rect 1900 5356 1908 5364
rect 1964 5356 1972 5364
rect 2236 5356 2244 5364
rect 2364 5356 2372 5364
rect 2588 5356 2596 5364
rect 2812 5356 2820 5364
rect 3100 5356 3108 5364
rect 3356 5356 3364 5364
rect 3740 5356 3748 5364
rect 3804 5356 3812 5364
rect 3948 5356 3956 5364
rect 4188 5356 4196 5364
rect 4284 5356 4292 5364
rect 28 5336 36 5344
rect 60 5336 68 5344
rect 156 5336 164 5344
rect 332 5336 340 5344
rect 428 5336 436 5344
rect 476 5336 484 5344
rect 524 5336 532 5344
rect 620 5336 628 5344
rect 732 5336 740 5344
rect 828 5336 836 5344
rect 844 5336 852 5344
rect 924 5336 932 5344
rect 1036 5336 1044 5344
rect 1132 5336 1140 5344
rect 1196 5336 1204 5344
rect 1212 5336 1220 5344
rect 1292 5336 1300 5344
rect 1308 5336 1316 5344
rect 1356 5336 1364 5344
rect 1420 5336 1428 5344
rect 1516 5336 1524 5344
rect 1692 5336 1700 5344
rect 1868 5336 1876 5344
rect 1916 5336 1924 5344
rect 2044 5336 2052 5344
rect 2204 5336 2212 5344
rect 2332 5336 2340 5344
rect 2444 5336 2452 5344
rect 2508 5336 2516 5344
rect 2620 5336 2628 5344
rect 2844 5336 2852 5344
rect 3004 5336 3012 5344
rect 3228 5336 3236 5344
rect 3340 5336 3348 5344
rect 3420 5336 3428 5344
rect 3516 5336 3524 5344
rect 12 5316 20 5324
rect 44 5316 52 5324
rect 92 5316 100 5324
rect 172 5316 180 5324
rect 316 5316 324 5324
rect 396 5316 404 5324
rect 540 5316 548 5324
rect 556 5316 564 5324
rect 892 5316 900 5324
rect 1068 5316 1076 5324
rect 1116 5316 1124 5324
rect 1180 5316 1188 5324
rect 3644 5336 3652 5344
rect 3692 5336 3700 5344
rect 3772 5336 3780 5344
rect 3788 5336 3796 5344
rect 3884 5336 3892 5344
rect 3980 5336 3988 5344
rect 4156 5336 4164 5344
rect 4204 5336 4212 5344
rect 4284 5336 4292 5344
rect 4300 5336 4308 5344
rect 4412 5336 4420 5344
rect 4460 5356 4468 5364
rect 4604 5356 4612 5364
rect 4892 5356 4900 5364
rect 5036 5356 5044 5364
rect 5212 5356 5220 5364
rect 5356 5356 5364 5364
rect 5740 5356 5748 5364
rect 5852 5356 5860 5364
rect 6044 5356 6052 5364
rect 4572 5336 4580 5344
rect 4732 5336 4740 5344
rect 4844 5336 4852 5344
rect 4860 5336 4868 5344
rect 4892 5336 4900 5344
rect 4908 5336 4916 5344
rect 4972 5336 4980 5344
rect 5068 5336 5076 5344
rect 5180 5336 5188 5344
rect 5228 5336 5236 5344
rect 5292 5336 5300 5344
rect 5340 5336 5348 5344
rect 5420 5336 5428 5344
rect 5468 5336 5476 5344
rect 5548 5336 5556 5344
rect 5580 5336 5588 5344
rect 5708 5336 5716 5344
rect 5820 5336 5828 5344
rect 5884 5336 5892 5344
rect 5916 5336 5924 5344
rect 5948 5336 5956 5344
rect 6012 5336 6020 5344
rect 6220 5336 6228 5344
rect 1308 5316 1316 5324
rect 1420 5316 1428 5324
rect 1436 5316 1444 5324
rect 1484 5316 1492 5324
rect 1564 5316 1572 5324
rect 1644 5316 1652 5324
rect 1692 5316 1700 5324
rect 1740 5316 1748 5324
rect 1820 5316 1828 5324
rect 1852 5316 1860 5324
rect 2012 5316 2020 5324
rect 2092 5316 2100 5324
rect 2140 5316 2148 5324
rect 2188 5316 2196 5324
rect 2268 5316 2276 5324
rect 2316 5316 2324 5324
rect 2364 5316 2372 5324
rect 2396 5316 2404 5324
rect 2556 5316 2564 5324
rect 2652 5316 2660 5324
rect 2700 5316 2708 5324
rect 2780 5316 2788 5324
rect 2860 5316 2868 5324
rect 2892 5316 2900 5324
rect 2956 5316 2964 5324
rect 3020 5316 3028 5324
rect 3068 5316 3076 5324
rect 3180 5316 3188 5324
rect 3212 5316 3220 5324
rect 3276 5316 3284 5324
rect 3628 5316 3636 5324
rect 3676 5316 3684 5324
rect 3708 5316 3716 5324
rect 3740 5316 3748 5324
rect 3836 5316 3844 5324
rect 3900 5316 3908 5324
rect 3996 5316 4004 5324
rect 4108 5316 4116 5324
rect 4140 5316 4148 5324
rect 4220 5316 4228 5324
rect 396 5296 404 5304
rect 444 5296 452 5304
rect 492 5296 500 5304
rect 572 5296 580 5304
rect 1084 5296 1092 5304
rect 1148 5296 1156 5304
rect 1244 5296 1252 5304
rect 1340 5296 1348 5304
rect 1404 5296 1412 5304
rect 1468 5296 1476 5304
rect 1596 5296 1604 5304
rect 1724 5296 1732 5304
rect 1836 5296 1844 5304
rect 1948 5296 1956 5304
rect 1980 5296 1988 5304
rect 1996 5296 2004 5304
rect 2108 5296 2116 5304
rect 2172 5296 2180 5304
rect 2252 5296 2260 5304
rect 2380 5296 2388 5304
rect 2476 5296 2484 5304
rect 2668 5296 2676 5304
rect 2684 5296 2692 5304
rect 2796 5296 2804 5304
rect 2876 5296 2884 5304
rect 2940 5296 2948 5304
rect 3052 5296 3060 5304
rect 3292 5296 3300 5304
rect 3308 5296 3316 5304
rect 3404 5296 3412 5304
rect 3484 5296 3492 5304
rect 3676 5296 3684 5304
rect 3740 5296 3748 5304
rect 3820 5296 3828 5304
rect 3868 5296 3876 5304
rect 3932 5296 3940 5304
rect 4124 5296 4132 5304
rect 4316 5316 4324 5324
rect 4380 5316 4388 5324
rect 4476 5316 4484 5324
rect 4508 5316 4516 5324
rect 4556 5316 4564 5324
rect 4684 5316 4692 5324
rect 4828 5316 4836 5324
rect 4924 5316 4932 5324
rect 4972 5316 4980 5324
rect 5084 5316 5092 5324
rect 5116 5316 5124 5324
rect 5164 5316 5172 5324
rect 5228 5316 5236 5324
rect 5308 5316 5316 5324
rect 5436 5316 5444 5324
rect 5484 5316 5492 5324
rect 5548 5316 5556 5324
rect 5644 5316 5652 5324
rect 5692 5316 5700 5324
rect 5788 5316 5796 5324
rect 5948 5316 5956 5324
rect 6044 5318 6052 5326
rect 4492 5296 4500 5304
rect 4620 5296 4628 5304
rect 4956 5296 4964 5304
rect 5020 5296 5028 5304
rect 5100 5296 5108 5304
rect 5276 5296 5284 5304
rect 5340 5296 5348 5304
rect 5500 5296 5508 5304
rect 5564 5296 5572 5304
rect 5612 5296 5620 5304
rect 5676 5296 5684 5304
rect 5804 5296 5812 5304
rect 5852 5296 5860 5304
rect 5980 5296 5988 5304
rect 6188 5296 6196 5304
rect 220 5276 228 5284
rect 1516 5276 1524 5284
rect 1660 5276 1668 5284
rect 1756 5276 1764 5284
rect 1772 5276 1780 5284
rect 1804 5276 1812 5284
rect 1916 5276 1924 5284
rect 2028 5276 2036 5284
rect 2076 5276 2084 5284
rect 2156 5276 2164 5284
rect 2284 5276 2292 5284
rect 2412 5276 2420 5284
rect 2716 5276 2724 5284
rect 2764 5276 2772 5284
rect 2908 5276 2916 5284
rect 2972 5276 2980 5284
rect 3260 5276 3268 5284
rect 3324 5276 3332 5284
rect 3852 5276 3860 5284
rect 4092 5276 4100 5284
rect 4524 5276 4532 5284
rect 4700 5276 4708 5284
rect 5132 5276 5140 5284
rect 5468 5276 5476 5284
rect 5532 5276 5540 5284
rect 5660 5276 5668 5284
rect 5772 5276 5780 5284
rect 1820 5256 1828 5264
rect 5820 5276 5828 5284
rect 1052 5236 1060 5244
rect 2732 5236 2740 5244
rect 2780 5236 2788 5244
rect 2892 5236 2900 5244
rect 2988 5236 2996 5244
rect 3180 5236 3188 5244
rect 3244 5236 3252 5244
rect 4988 5236 4996 5244
rect 5148 5236 5156 5244
rect 5244 5236 5252 5244
rect 6204 5236 6212 5244
rect 1566 5206 1574 5214
rect 1580 5206 1588 5214
rect 1594 5206 1602 5214
rect 4638 5206 4646 5214
rect 4652 5206 4660 5214
rect 4666 5206 4674 5214
rect 28 5176 36 5184
rect 252 5176 260 5184
rect 284 5176 292 5184
rect 348 5176 356 5184
rect 412 5176 420 5184
rect 636 5176 644 5184
rect 1372 5176 1380 5184
rect 1692 5176 1700 5184
rect 1996 5176 2004 5184
rect 2076 5176 2084 5184
rect 2124 5176 2132 5184
rect 2172 5176 2180 5184
rect 2492 5176 2500 5184
rect 3500 5176 3508 5184
rect 3692 5176 3700 5184
rect 3756 5176 3764 5184
rect 3916 5176 3924 5184
rect 3964 5176 3972 5184
rect 4268 5176 4276 5184
rect 4716 5176 4724 5184
rect 4796 5176 4804 5184
rect 4828 5176 4836 5184
rect 4892 5176 4900 5184
rect 5052 5176 5060 5184
rect 5340 5176 5348 5184
rect 5468 5176 5476 5184
rect 5660 5176 5668 5184
rect 5756 5176 5764 5184
rect 5772 5176 5780 5184
rect 5852 5176 5860 5184
rect 6012 5176 6020 5184
rect 6220 5176 6228 5184
rect 3868 5156 3876 5164
rect 4476 5156 4484 5164
rect 4540 5156 4548 5164
rect 828 5136 836 5144
rect 924 5136 932 5144
rect 3324 5136 3332 5144
rect 3436 5136 3444 5144
rect 3484 5136 3492 5144
rect 3740 5136 3748 5144
rect 3852 5136 3860 5144
rect 4252 5136 4260 5144
rect 4300 5136 4308 5144
rect 4460 5136 4468 5144
rect 4524 5136 4532 5144
rect 4700 5136 4708 5144
rect 4844 5136 4852 5144
rect 4908 5136 4916 5144
rect 5036 5136 5044 5144
rect 5452 5136 5460 5144
rect 5516 5136 5524 5144
rect 5548 5136 5556 5144
rect 5676 5136 5684 5144
rect 5740 5136 5748 5144
rect 6236 5136 6244 5144
rect 220 5116 228 5124
rect 332 5116 340 5124
rect 588 5116 596 5124
rect 716 5116 724 5124
rect 892 5116 900 5124
rect 956 5116 964 5124
rect 988 5116 996 5124
rect 60 5096 68 5104
rect 220 5096 228 5104
rect 252 5096 260 5104
rect 284 5096 292 5104
rect 380 5096 388 5104
rect 428 5096 436 5104
rect 460 5096 468 5104
rect 476 5096 484 5104
rect 492 5096 500 5104
rect 828 5096 836 5104
rect 860 5096 868 5104
rect 956 5096 964 5104
rect 1068 5116 1076 5124
rect 1132 5116 1140 5124
rect 1196 5116 1204 5124
rect 1244 5116 1252 5124
rect 1340 5116 1348 5124
rect 1052 5096 1060 5104
rect 1100 5096 1108 5104
rect 1148 5096 1156 5104
rect 1164 5096 1172 5104
rect 1180 5096 1188 5104
rect 1308 5096 1316 5104
rect 1324 5096 1332 5104
rect 1372 5096 1380 5104
rect 1468 5116 1476 5124
rect 1836 5116 1844 5124
rect 1916 5116 1924 5124
rect 1948 5116 1956 5124
rect 2060 5116 2068 5124
rect 2140 5116 2148 5124
rect 2204 5116 2212 5124
rect 2284 5116 2292 5124
rect 2524 5116 2532 5124
rect 2620 5116 2628 5124
rect 3052 5116 3060 5124
rect 3244 5116 3252 5124
rect 3260 5116 3268 5124
rect 3356 5116 3364 5124
rect 3372 5116 3380 5124
rect 3452 5116 3460 5124
rect 3516 5116 3524 5124
rect 3628 5116 3636 5124
rect 3708 5116 3716 5124
rect 3884 5116 3892 5124
rect 3932 5116 3940 5124
rect 4060 5116 4068 5124
rect 4076 5116 4084 5124
rect 4140 5116 4148 5124
rect 4204 5116 4212 5124
rect 4220 5116 4228 5124
rect 4332 5116 4340 5124
rect 4396 5116 4404 5124
rect 4428 5116 4436 5124
rect 4492 5116 4500 5124
rect 4556 5116 4564 5124
rect 4732 5116 4740 5124
rect 4812 5116 4820 5124
rect 4876 5116 4884 5124
rect 5004 5116 5012 5124
rect 5212 5116 5220 5124
rect 5420 5116 5428 5124
rect 5484 5116 5492 5124
rect 5612 5116 5620 5124
rect 5628 5116 5636 5124
rect 5708 5116 5716 5124
rect 5868 5116 5876 5124
rect 5932 5116 5940 5124
rect 6204 5116 6212 5124
rect 1420 5096 1428 5104
rect 1676 5096 1684 5104
rect 1740 5096 1748 5104
rect 1756 5096 1764 5104
rect 1820 5096 1828 5104
rect 1964 5096 1972 5104
rect 1996 5096 2004 5104
rect 2188 5096 2196 5104
rect 2316 5096 2324 5104
rect 2412 5096 2420 5104
rect 2444 5096 2452 5104
rect 2588 5096 2596 5104
rect 2684 5096 2692 5104
rect 2828 5096 2836 5104
rect 2972 5096 2980 5104
rect 3036 5096 3044 5104
rect 3164 5096 3172 5104
rect 3260 5096 3268 5104
rect 3340 5096 3348 5104
rect 12 5076 20 5084
rect 76 5076 84 5084
rect 204 5076 212 5084
rect 268 5076 276 5084
rect 364 5076 372 5084
rect 380 5076 388 5084
rect 444 5076 452 5084
rect 492 5076 500 5084
rect 556 5076 564 5084
rect 604 5076 612 5084
rect 700 5076 708 5084
rect 748 5076 756 5084
rect 780 5076 788 5084
rect 892 5076 900 5084
rect 924 5076 932 5084
rect 940 5076 948 5084
rect 1004 5076 1012 5084
rect 1052 5076 1060 5084
rect 1068 5076 1076 5084
rect 1116 5076 1124 5084
rect 1180 5076 1188 5084
rect 1228 5076 1236 5084
rect 1276 5076 1284 5084
rect 1292 5076 1300 5084
rect 1356 5076 1364 5084
rect 1420 5076 1428 5084
rect 1580 5076 1588 5084
rect 1724 5076 1732 5084
rect 1804 5076 1812 5084
rect 1868 5076 1876 5084
rect 1916 5076 1924 5084
rect 2060 5076 2068 5084
rect 2092 5076 2100 5084
rect 2188 5076 2196 5084
rect 2236 5076 2244 5084
rect 2364 5076 2372 5084
rect 2444 5076 2452 5084
rect 92 5056 100 5064
rect 316 5056 324 5064
rect 508 5056 516 5064
rect 540 5056 548 5064
rect 732 5056 740 5064
rect 764 5056 772 5064
rect 1644 5056 1652 5064
rect 1788 5056 1796 5064
rect 1852 5056 1860 5064
rect 2044 5056 2052 5064
rect 2268 5056 2276 5064
rect 2428 5056 2436 5064
rect 2572 5076 2580 5084
rect 2604 5076 2612 5084
rect 2668 5076 2676 5084
rect 2796 5076 2804 5084
rect 2540 5056 2548 5064
rect 2652 5056 2660 5064
rect 2764 5056 2772 5064
rect 2908 5056 2916 5064
rect 2956 5076 2964 5084
rect 2972 5076 2980 5084
rect 3020 5076 3028 5084
rect 3084 5076 3092 5084
rect 3148 5076 3156 5084
rect 3212 5076 3220 5084
rect 3244 5076 3252 5084
rect 3292 5076 3300 5084
rect 3340 5076 3348 5084
rect 3420 5096 3428 5104
rect 3500 5096 3508 5104
rect 3548 5096 3556 5104
rect 3580 5096 3588 5104
rect 3644 5096 3652 5104
rect 3724 5096 3732 5104
rect 3772 5096 3780 5104
rect 3868 5096 3876 5104
rect 3964 5096 3972 5104
rect 4108 5096 4116 5104
rect 4156 5096 4164 5104
rect 4236 5096 4244 5104
rect 4300 5096 4308 5104
rect 4364 5096 4372 5104
rect 4476 5096 4484 5104
rect 4540 5096 4548 5104
rect 4620 5096 4628 5104
rect 4716 5096 4724 5104
rect 4748 5096 4756 5104
rect 4828 5096 4836 5104
rect 4892 5096 4900 5104
rect 4940 5096 4948 5104
rect 4972 5096 4980 5104
rect 5020 5096 5028 5104
rect 5436 5096 5444 5104
rect 5500 5096 5508 5104
rect 5532 5096 5540 5104
rect 5660 5096 5668 5104
rect 5724 5096 5732 5104
rect 5804 5096 5812 5104
rect 5900 5096 5908 5104
rect 5980 5096 5988 5104
rect 6220 5096 6228 5104
rect 3420 5076 3428 5084
rect 3564 5076 3572 5084
rect 3644 5076 3652 5084
rect 3660 5076 3668 5084
rect 3788 5076 3796 5084
rect 3820 5076 3828 5084
rect 3980 5076 3988 5084
rect 3996 5076 4004 5084
rect 4044 5076 4052 5084
rect 4092 5076 4100 5084
rect 4172 5076 4180 5084
rect 4284 5076 4292 5084
rect 4348 5076 4356 5084
rect 4380 5076 4388 5084
rect 4588 5076 4596 5084
rect 4604 5076 4612 5084
rect 4764 5076 4772 5084
rect 4956 5076 4964 5084
rect 5068 5076 5076 5084
rect 5404 5076 5412 5084
rect 5580 5080 5588 5088
rect 5596 5076 5604 5084
rect 5820 5076 5828 5084
rect 5836 5076 5844 5084
rect 5868 5076 5876 5084
rect 5948 5076 5956 5084
rect 6044 5076 6052 5084
rect 6092 5076 6100 5084
rect 6188 5076 6196 5084
rect 2988 5056 2996 5064
rect 3372 5056 3380 5064
rect 3532 5056 3540 5064
rect 3692 5056 3700 5064
rect 3820 5056 3828 5064
rect 3900 5056 3908 5064
rect 4060 5056 4068 5064
rect 4204 5056 4212 5064
rect 4428 5056 4436 5064
rect 4572 5056 4580 5064
rect 4796 5056 4804 5064
rect 4988 5056 4996 5064
rect 5196 5056 5204 5064
rect 5260 5056 5268 5064
rect 5292 5056 5300 5064
rect 5628 5056 5636 5064
rect 6076 5056 6084 5064
rect 572 5036 580 5044
rect 1244 5036 1252 5044
rect 1516 5036 1524 5044
rect 2252 5036 2260 5044
rect 2284 5036 2292 5044
rect 2428 5036 2436 5044
rect 2556 5036 2564 5044
rect 2668 5036 2676 5044
rect 2780 5036 2788 5044
rect 2860 5036 2868 5044
rect 2940 5036 2948 5044
rect 3052 5036 3060 5044
rect 3196 5036 3204 5044
rect 5132 5036 5140 5044
rect 6060 5036 6068 5044
rect 6124 5036 6132 5044
rect 3118 5006 3126 5014
rect 3132 5006 3140 5014
rect 3146 5006 3154 5014
rect 60 4976 68 4984
rect 124 4976 132 4984
rect 188 4976 196 4984
rect 332 4976 340 4984
rect 396 4976 404 4984
rect 444 4976 452 4984
rect 460 4976 468 4984
rect 540 4976 548 4984
rect 604 4976 612 4984
rect 892 4976 900 4984
rect 956 4976 964 4984
rect 1052 4976 1060 4984
rect 1084 4976 1092 4984
rect 1596 4976 1604 4984
rect 1708 4976 1716 4984
rect 1772 4976 1780 4984
rect 1916 4976 1924 4984
rect 2172 4976 2180 4984
rect 2700 4976 2708 4984
rect 3116 4976 3124 4984
rect 3308 4976 3316 4984
rect 3500 4976 3508 4984
rect 3532 4976 3540 4984
rect 3676 4976 3684 4984
rect 3804 4976 3812 4984
rect 3852 4976 3860 4984
rect 4188 4976 4196 4984
rect 4284 4976 4292 4984
rect 4348 4976 4356 4984
rect 4604 4976 4612 4984
rect 4620 4976 4628 4984
rect 4716 4976 4724 4984
rect 4940 4976 4948 4984
rect 4988 4976 4996 4984
rect 5084 4976 5092 4984
rect 5148 4976 5156 4984
rect 5180 4976 5188 4984
rect 5212 4976 5220 4984
rect 5340 4976 5348 4984
rect 5516 4976 5524 4984
rect 5580 4976 5588 4984
rect 5804 4976 5812 4984
rect 5868 4976 5876 4984
rect 5980 4976 5988 4984
rect 6044 4976 6052 4984
rect 6108 4976 6116 4984
rect 204 4956 212 4964
rect 412 4956 420 4964
rect 1036 4956 1044 4964
rect 1068 4956 1076 4964
rect 1164 4956 1172 4964
rect 1372 4956 1380 4964
rect 1580 4956 1588 4964
rect 1836 4956 1844 4964
rect 1932 4956 1940 4964
rect 2188 4956 2196 4964
rect 2236 4956 2244 4964
rect 2380 4956 2388 4964
rect 2524 4956 2532 4964
rect 2860 4956 2868 4964
rect 3580 4956 3588 4964
rect 3612 4956 3620 4964
rect 3820 4956 3828 4964
rect 3916 4956 3924 4964
rect 3996 4956 4004 4964
rect 4300 4956 4308 4964
rect 4364 4956 4372 4964
rect 4444 4956 4452 4964
rect 4540 4956 4548 4964
rect 4652 4956 4660 4964
rect 12 4936 20 4944
rect 108 4936 116 4944
rect 156 4936 164 4944
rect 220 4936 228 4944
rect 316 4936 324 4944
rect 364 4936 372 4944
rect 508 4936 516 4944
rect 524 4936 532 4944
rect 572 4936 580 4944
rect 668 4936 676 4944
rect 716 4936 724 4944
rect 732 4936 740 4944
rect 172 4916 180 4924
rect 380 4916 388 4924
rect 492 4916 500 4924
rect 844 4936 852 4944
rect 924 4936 932 4944
rect 972 4936 980 4944
rect 988 4936 996 4944
rect 1100 4936 1108 4944
rect 1148 4936 1156 4944
rect 1244 4936 1252 4944
rect 1308 4936 1316 4944
rect 1436 4936 1444 4944
rect 1468 4936 1476 4944
rect 1484 4936 1492 4944
rect 1548 4936 1556 4944
rect 1724 4936 1732 4944
rect 1820 4936 1828 4944
rect 1868 4936 1876 4944
rect 1964 4936 1972 4944
rect 2092 4936 2100 4944
rect 2156 4936 2164 4944
rect 2348 4936 2356 4944
rect 2380 4936 2388 4944
rect 2572 4936 2580 4944
rect 2636 4936 2644 4944
rect 2652 4936 2660 4944
rect 2732 4936 2740 4944
rect 2780 4936 2788 4944
rect 2924 4936 2932 4944
rect 2988 4936 2996 4944
rect 3004 4936 3012 4944
rect 3052 4936 3060 4944
rect 3180 4936 3188 4944
rect 3276 4936 3284 4944
rect 3372 4936 3380 4944
rect 3404 4936 3412 4944
rect 3452 4936 3460 4944
rect 3788 4936 3796 4944
rect 3852 4936 3860 4944
rect 3884 4936 3892 4944
rect 3916 4936 3924 4944
rect 3948 4936 3956 4944
rect 3980 4936 3988 4944
rect 4012 4936 4020 4944
rect 4060 4936 4068 4944
rect 4092 4936 4100 4944
rect 4156 4936 4164 4944
rect 4204 4936 4212 4944
rect 4220 4936 4228 4944
rect 4332 4936 4340 4944
rect 4460 4936 4468 4944
rect 4572 4936 4580 4944
rect 4636 4936 4644 4944
rect 4732 4936 4740 4944
rect 4780 4956 4788 4964
rect 4924 4956 4932 4964
rect 5356 4956 5364 4964
rect 5612 4956 5620 4964
rect 5884 4956 5892 4964
rect 1212 4916 1220 4924
rect 1260 4916 1268 4924
rect 1324 4916 1332 4924
rect 1404 4916 1412 4924
rect 1452 4916 1460 4924
rect 1484 4916 1492 4924
rect 1628 4916 1636 4924
rect 1884 4916 1892 4924
rect 1964 4916 1972 4924
rect 1980 4916 1988 4924
rect 2060 4916 2068 4924
rect 2140 4916 2148 4924
rect 2236 4916 2244 4924
rect 2300 4916 2308 4924
rect 2332 4916 2340 4924
rect 2428 4916 2436 4924
rect 2492 4916 2500 4924
rect 2572 4916 2580 4924
rect 2620 4916 2628 4924
rect 4860 4936 4868 4944
rect 4956 4936 4964 4944
rect 5020 4936 5028 4944
rect 5036 4936 5044 4944
rect 5100 4936 5108 4944
rect 5164 4936 5172 4944
rect 5324 4936 5332 4944
rect 5420 4936 5428 4944
rect 5500 4936 5508 4944
rect 5852 4936 5860 4944
rect 6028 4936 6036 4944
rect 6172 4936 6180 4944
rect 2796 4916 2804 4924
rect 2812 4916 2820 4924
rect 2908 4916 2916 4924
rect 2972 4916 2980 4924
rect 3228 4916 3236 4924
rect 3420 4916 3428 4924
rect 3468 4916 3476 4924
rect 3532 4916 3540 4924
rect 3580 4916 3588 4924
rect 3660 4916 3668 4924
rect 3724 4916 3732 4924
rect 3772 4916 3780 4924
rect 3836 4916 3844 4924
rect 3900 4916 3908 4924
rect 3964 4916 3972 4924
rect 4028 4916 4036 4924
rect 4076 4916 4084 4924
rect 4092 4916 4100 4924
rect 4140 4916 4148 4924
rect 4236 4916 4244 4924
rect 4252 4916 4260 4924
rect 4316 4916 4324 4924
rect 4412 4916 4420 4924
rect 4540 4916 4548 4924
rect 4780 4916 4788 4924
rect 4812 4916 4820 4924
rect 4972 4916 4980 4924
rect 5052 4916 5060 4924
rect 5116 4916 5124 4924
rect 5292 4916 5300 4924
rect 5388 4916 5396 4924
rect 5452 4916 5460 4924
rect 5580 4916 5588 4924
rect 5612 4916 5620 4924
rect 5660 4916 5668 4924
rect 5740 4916 5748 4924
rect 5804 4916 5812 4924
rect 5836 4916 5844 4924
rect 5932 4916 5940 4924
rect 5964 4916 5972 4924
rect 5980 4916 5988 4924
rect 6204 4916 6212 4924
rect 124 4896 132 4904
rect 332 4896 340 4904
rect 556 4896 564 4904
rect 684 4896 692 4904
rect 700 4896 708 4904
rect 892 4896 900 4904
rect 940 4896 948 4904
rect 1020 4896 1028 4904
rect 1036 4896 1044 4904
rect 1148 4896 1156 4904
rect 1356 4896 1364 4904
rect 1420 4896 1428 4904
rect 1532 4896 1540 4904
rect 1580 4896 1588 4904
rect 1916 4896 1924 4904
rect 2012 4896 2020 4904
rect 2076 4896 2084 4904
rect 2108 4896 2116 4904
rect 2124 4896 2132 4904
rect 2252 4896 2260 4904
rect 2316 4896 2324 4904
rect 2444 4896 2452 4904
rect 2508 4896 2516 4904
rect 2524 4896 2532 4904
rect 2588 4896 2596 4904
rect 2700 4896 2708 4904
rect 2716 4896 2724 4904
rect 2844 4896 2852 4904
rect 2876 4896 2884 4904
rect 2940 4896 2948 4904
rect 2972 4896 2980 4904
rect 3036 4896 3044 4904
rect 3212 4896 3220 4904
rect 3436 4896 3444 4904
rect 3500 4896 3508 4904
rect 3516 4896 3524 4904
rect 3644 4896 3652 4904
rect 3708 4896 3716 4904
rect 3916 4896 3924 4904
rect 4044 4896 4052 4904
rect 4156 4896 4164 4904
rect 4268 4896 4276 4904
rect 4428 4896 4436 4904
rect 4556 4896 4564 4904
rect 4604 4896 4612 4904
rect 4700 4896 4708 4904
rect 4908 4896 4916 4904
rect 4988 4896 4996 4904
rect 5148 4896 5156 4904
rect 5196 4896 5204 4904
rect 5212 4896 5220 4904
rect 5244 4896 5252 4904
rect 5372 4896 5380 4904
rect 5436 4896 5444 4904
rect 5596 4896 5604 4904
rect 5692 4896 5700 4904
rect 5740 4896 5748 4904
rect 5804 4896 5812 4904
rect 5932 4896 5940 4904
rect 284 4876 292 4884
rect 764 4876 772 4884
rect 2028 4876 2036 4884
rect 2060 4876 2068 4884
rect 2092 4876 2100 4884
rect 2220 4876 2228 4884
rect 2284 4876 2292 4884
rect 2412 4876 2420 4884
rect 2476 4876 2484 4884
rect 3196 4876 3204 4884
rect 3404 4876 3412 4884
rect 3548 4876 3556 4884
rect 3644 4876 3652 4884
rect 3676 4876 3684 4884
rect 3740 4876 3748 4884
rect 4396 4876 4404 4884
rect 4492 4876 4500 4884
rect 4524 4876 4532 4884
rect 4876 4876 4884 4884
rect 5404 4876 5412 4884
rect 5468 4876 5476 4884
rect 5564 4876 5572 4884
rect 5644 4876 5652 4884
rect 5724 4876 5732 4884
rect 5788 4876 5796 4884
rect 5916 4876 5924 4884
rect 6060 4896 6068 4904
rect 6188 4896 6196 4904
rect 2300 4856 2308 4864
rect 4412 4856 4420 4864
rect 5996 4876 6004 4884
rect 6220 4876 6228 4884
rect 1292 4836 1300 4844
rect 1324 4836 1332 4844
rect 1404 4836 1412 4844
rect 1980 4836 1988 4844
rect 2428 4836 2436 4844
rect 2492 4836 2500 4844
rect 2620 4836 2628 4844
rect 2908 4836 2916 4844
rect 3020 4836 3028 4844
rect 3260 4836 3268 4844
rect 5484 4836 5492 4844
rect 5740 4836 5748 4844
rect 5804 4836 5812 4844
rect 6204 4836 6212 4844
rect 1566 4806 1574 4814
rect 1580 4806 1588 4814
rect 1594 4806 1602 4814
rect 4638 4806 4646 4814
rect 4652 4806 4660 4814
rect 4666 4806 4674 4814
rect 76 4776 84 4784
rect 492 4776 500 4784
rect 748 4776 756 4784
rect 1084 4776 1092 4784
rect 1372 4776 1380 4784
rect 1500 4776 1508 4784
rect 1852 4776 1860 4784
rect 1932 4776 1940 4784
rect 1980 4776 1988 4784
rect 2060 4776 2068 4784
rect 2524 4776 2532 4784
rect 3036 4776 3044 4784
rect 3228 4776 3236 4784
rect 3468 4776 3476 4784
rect 3500 4776 3508 4784
rect 3564 4776 3572 4784
rect 3644 4776 3652 4784
rect 4316 4776 4324 4784
rect 4572 4776 4580 4784
rect 4828 4776 4836 4784
rect 4940 4776 4948 4784
rect 5084 4776 5092 4784
rect 5148 4776 5156 4784
rect 5436 4776 5444 4784
rect 5628 4776 5636 4784
rect 5852 4776 5860 4784
rect 5932 4776 5940 4784
rect 6140 4776 6148 4784
rect 2652 4756 2660 4764
rect 3772 4756 3780 4764
rect 4060 4756 4068 4764
rect 4252 4756 4260 4764
rect 4380 4756 4388 4764
rect 476 4736 484 4744
rect 636 4736 644 4744
rect 940 4736 948 4744
rect 1004 4736 1012 4744
rect 1420 4736 1428 4744
rect 1516 4736 1524 4744
rect 1772 4736 1780 4744
rect 1836 4736 1844 4744
rect 1964 4736 1972 4744
rect 2012 4736 2020 4744
rect 2044 4736 2052 4744
rect 2124 4736 2132 4744
rect 2460 4736 2468 4744
rect 2508 4736 2516 4744
rect 2588 4736 2596 4744
rect 2636 4736 2644 4744
rect 2700 4736 2708 4744
rect 3020 4736 3028 4744
rect 3212 4736 3220 4744
rect 3356 4736 3364 4744
rect 3452 4736 3460 4744
rect 3628 4736 3636 4744
rect 3756 4736 3764 4744
rect 3820 4736 3828 4744
rect 3836 4736 3844 4744
rect 4044 4736 4052 4744
rect 4236 4736 4244 4744
rect 4300 4736 4308 4744
rect 4364 4736 4372 4744
rect 4556 4736 4564 4744
rect 4812 4736 4820 4744
rect 5068 4736 5076 4744
rect 5244 4736 5252 4744
rect 5836 4736 5844 4744
rect 5948 4736 5956 4744
rect 508 4716 516 4724
rect 524 4716 532 4724
rect 972 4716 980 4724
rect 1292 4716 1300 4724
rect 1388 4716 1396 4724
rect 1436 4716 1444 4724
rect 1516 4716 1524 4724
rect 1804 4716 1812 4724
rect 1868 4716 1876 4724
rect 1996 4716 2004 4724
rect 2092 4716 2100 4724
rect 2156 4716 2164 4724
rect 2204 4716 2212 4724
rect 2252 4716 2260 4724
rect 2476 4716 2484 4724
rect 2540 4716 2548 4724
rect 2556 4716 2564 4724
rect 2668 4716 2676 4724
rect 2732 4716 2740 4724
rect 2844 4716 2852 4724
rect 2988 4716 2996 4724
rect 3052 4716 3060 4724
rect 3244 4716 3252 4724
rect 3340 4716 3348 4724
rect 3420 4716 3428 4724
rect 3532 4716 3540 4724
rect 3596 4716 3604 4724
rect 3660 4716 3668 4724
rect 3788 4716 3796 4724
rect 3852 4716 3860 4724
rect 4012 4716 4020 4724
rect 4076 4716 4084 4724
rect 4204 4716 4212 4724
rect 4268 4716 4276 4724
rect 4332 4716 4340 4724
rect 4396 4716 4404 4724
rect 4460 4716 4468 4724
rect 4524 4716 4532 4724
rect 4588 4716 4596 4724
rect 4764 4716 4772 4724
rect 4780 4716 4788 4724
rect 5100 4716 5108 4724
rect 5276 4716 5284 4724
rect 5340 4716 5348 4724
rect 5740 4716 5748 4724
rect 5804 4716 5812 4724
rect 5900 4716 5908 4724
rect 5980 4716 5988 4724
rect 6108 4716 6116 4724
rect 188 4696 196 4704
rect 332 4696 340 4704
rect 492 4696 500 4704
rect 12 4676 20 4684
rect 108 4676 116 4684
rect 156 4680 164 4688
rect 188 4656 196 4664
rect 236 4676 244 4684
rect 348 4676 356 4684
rect 444 4676 452 4684
rect 556 4676 564 4684
rect 940 4696 948 4704
rect 972 4696 980 4704
rect 1084 4696 1092 4704
rect 1164 4696 1172 4704
rect 1308 4696 1316 4704
rect 1324 4696 1332 4704
rect 1404 4696 1412 4704
rect 1452 4696 1460 4704
rect 1532 4696 1540 4704
rect 1644 4696 1652 4704
rect 1676 4696 1684 4704
rect 1772 4696 1780 4704
rect 1852 4696 1860 4704
rect 1884 4696 1892 4704
rect 1980 4696 1988 4704
rect 2028 4696 2036 4704
rect 2140 4696 2148 4704
rect 2332 4696 2340 4704
rect 2460 4696 2468 4704
rect 2524 4696 2532 4704
rect 2572 4696 2580 4704
rect 2604 4696 2612 4704
rect 2652 4696 2660 4704
rect 2716 4696 2724 4704
rect 2748 4696 2756 4704
rect 2796 4696 2804 4704
rect 2956 4696 2964 4704
rect 3004 4696 3012 4704
rect 3084 4696 3092 4704
rect 3228 4696 3236 4704
rect 3260 4696 3268 4704
rect 3404 4696 3412 4704
rect 3436 4696 3444 4704
rect 3500 4696 3508 4704
rect 3564 4696 3572 4704
rect 3644 4696 3652 4704
rect 3676 4696 3684 4704
rect 3724 4696 3732 4704
rect 3772 4696 3780 4704
rect 3836 4696 3844 4704
rect 3932 4696 3940 4704
rect 4012 4696 4020 4704
rect 4060 4696 4068 4704
rect 4124 4696 4132 4704
rect 4252 4696 4260 4704
rect 4316 4696 4324 4704
rect 4380 4696 4388 4704
rect 4412 4696 4420 4704
rect 4476 4696 4484 4704
rect 4492 4696 4500 4704
rect 4572 4696 4580 4704
rect 4604 4696 4612 4704
rect 4636 4696 4644 4704
rect 4748 4696 4756 4704
rect 4796 4696 4804 4704
rect 4844 4696 4852 4704
rect 4908 4696 4916 4704
rect 5084 4696 5092 4704
rect 5244 4696 5252 4704
rect 5308 4696 5316 4704
rect 5420 4696 5428 4704
rect 5468 4696 5476 4704
rect 5500 4696 5508 4704
rect 5532 4696 5540 4704
rect 5548 4696 5556 4704
rect 5708 4696 5716 4704
rect 5756 4696 5764 4704
rect 5772 4696 5780 4704
rect 5788 4696 5796 4704
rect 5852 4696 5860 4704
rect 5932 4696 5940 4704
rect 6012 4696 6020 4704
rect 6044 4696 6052 4704
rect 6140 4696 6148 4704
rect 6156 4696 6164 4704
rect 6220 4696 6228 4704
rect 668 4676 676 4684
rect 684 4676 692 4684
rect 780 4676 788 4684
rect 844 4676 852 4684
rect 892 4676 900 4684
rect 876 4656 884 4664
rect 1196 4676 1204 4684
rect 1276 4676 1284 4684
rect 1340 4676 1348 4684
rect 1660 4676 1668 4684
rect 1756 4676 1764 4684
rect 1900 4676 1908 4684
rect 2140 4676 2148 4684
rect 2172 4676 2180 4684
rect 2220 4676 2228 4684
rect 2364 4676 2372 4684
rect 2764 4676 2772 4684
rect 2812 4676 2820 4684
rect 2940 4676 2948 4684
rect 3068 4676 3076 4684
rect 3100 4676 3108 4684
rect 3276 4676 3284 4684
rect 3324 4676 3332 4684
rect 3404 4676 3412 4684
rect 3484 4676 3492 4684
rect 3548 4676 3556 4684
rect 3692 4676 3700 4684
rect 3948 4676 3956 4684
rect 4108 4676 4116 4684
rect 4140 4676 4148 4684
rect 4172 4676 4180 4684
rect 4204 4676 4212 4684
rect 4412 4676 4420 4684
rect 4476 4676 4484 4684
rect 4524 4676 4532 4684
rect 4620 4676 4628 4684
rect 4652 4676 4660 4684
rect 4732 4676 4740 4684
rect 4860 4676 4868 4684
rect 4876 4676 4884 4684
rect 4892 4676 4900 4684
rect 4988 4676 4996 4684
rect 5036 4676 5044 4684
rect 5116 4676 5124 4684
rect 5212 4676 5220 4684
rect 5228 4676 5236 4684
rect 5292 4676 5300 4684
rect 5356 4676 5364 4684
rect 5372 4676 5380 4684
rect 5484 4676 5492 4684
rect 5516 4676 5524 4684
rect 5564 4676 5572 4684
rect 5580 4676 5588 4684
rect 5612 4676 5620 4684
rect 5660 4676 5668 4684
rect 5692 4676 5700 4684
rect 5756 4676 5764 4684
rect 6028 4676 6036 4684
rect 6060 4676 6068 4684
rect 6092 4676 6100 4684
rect 6156 4676 6164 4684
rect 6204 4676 6212 4684
rect 1004 4656 1012 4664
rect 1020 4656 1028 4664
rect 1052 4656 1060 4664
rect 1164 4656 1172 4664
rect 1292 4656 1300 4664
rect 1372 4656 1380 4664
rect 1500 4656 1508 4664
rect 1644 4656 1652 4664
rect 1932 4656 1940 4664
rect 2076 4656 2084 4664
rect 2204 4656 2212 4664
rect 2348 4656 2356 4664
rect 2796 4656 2804 4664
rect 2828 4656 2836 4664
rect 2956 4656 2964 4664
rect 3180 4656 3188 4664
rect 3308 4656 3316 4664
rect 3724 4656 3732 4664
rect 3836 4656 3844 4664
rect 3884 4656 3892 4664
rect 4924 4656 4932 4664
rect 4972 4656 4980 4664
rect 5356 4656 5364 4664
rect 5676 4656 5684 4664
rect 5900 4656 5908 4664
rect 6092 4656 6100 4664
rect 6172 4656 6180 4664
rect 124 4636 132 4644
rect 268 4636 276 4644
rect 1036 4636 1044 4644
rect 1180 4636 1188 4644
rect 1660 4636 1668 4644
rect 2252 4636 2260 4644
rect 2300 4636 2308 4644
rect 2412 4636 2420 4644
rect 2460 4636 2468 4644
rect 2716 4636 2724 4644
rect 2892 4636 2900 4644
rect 3900 4636 3908 4644
rect 5020 4636 5028 4644
rect 5980 4636 5988 4644
rect 3118 4606 3126 4614
rect 3132 4606 3140 4614
rect 3146 4606 3154 4614
rect 76 4576 84 4584
rect 220 4576 228 4584
rect 268 4576 276 4584
rect 348 4576 356 4584
rect 444 4576 452 4584
rect 620 4576 628 4584
rect 828 4576 836 4584
rect 1020 4576 1028 4584
rect 1100 4576 1108 4584
rect 1132 4576 1140 4584
rect 1324 4576 1332 4584
rect 1436 4576 1444 4584
rect 1516 4576 1524 4584
rect 1612 4576 1620 4584
rect 1740 4576 1748 4584
rect 2140 4576 2148 4584
rect 2332 4576 2340 4584
rect 2636 4576 2644 4584
rect 2700 4576 2708 4584
rect 3436 4576 3444 4584
rect 3548 4576 3556 4584
rect 3612 4576 3620 4584
rect 3740 4576 3748 4584
rect 3852 4576 3860 4584
rect 3932 4576 3940 4584
rect 3964 4576 3972 4584
rect 4108 4576 4116 4584
rect 4172 4576 4180 4584
rect 4284 4576 4292 4584
rect 4380 4576 4388 4584
rect 4460 4576 4468 4584
rect 4508 4576 4516 4584
rect 4604 4576 4612 4584
rect 4732 4576 4740 4584
rect 4764 4576 4772 4584
rect 4828 4576 4836 4584
rect 4892 4576 4900 4584
rect 4924 4576 4932 4584
rect 4972 4576 4980 4584
rect 5068 4576 5076 4584
rect 5100 4576 5108 4584
rect 5164 4576 5172 4584
rect 5276 4576 5284 4584
rect 5340 4576 5348 4584
rect 5436 4576 5444 4584
rect 5580 4576 5588 4584
rect 5612 4576 5620 4584
rect 5660 4576 5668 4584
rect 5692 4576 5700 4584
rect 5900 4576 5908 4584
rect 5932 4576 5940 4584
rect 636 4556 644 4564
rect 1036 4556 1044 4564
rect 1116 4556 1124 4564
rect 1228 4556 1236 4564
rect 1324 4556 1332 4564
rect 12 4536 20 4544
rect 108 4536 116 4544
rect 124 4536 132 4544
rect 236 4536 244 4544
rect 284 4536 292 4544
rect 396 4536 404 4544
rect 604 4536 612 4544
rect 700 4536 708 4544
rect 748 4536 756 4544
rect 764 4536 772 4544
rect 860 4536 868 4544
rect 876 4536 884 4544
rect 972 4536 980 4544
rect 1004 4536 1012 4544
rect 1148 4536 1156 4544
rect 140 4516 148 4524
rect 412 4516 420 4524
rect 476 4516 484 4524
rect 556 4516 564 4524
rect 588 4516 596 4524
rect 684 4516 692 4524
rect 988 4516 996 4524
rect 1068 4516 1076 4524
rect 1164 4516 1172 4524
rect 1196 4536 1204 4544
rect 1260 4536 1268 4544
rect 1340 4536 1348 4544
rect 1596 4556 1604 4564
rect 1740 4556 1748 4564
rect 1420 4536 1428 4544
rect 1484 4536 1492 4544
rect 1532 4536 1540 4544
rect 1628 4536 1636 4544
rect 1756 4536 1764 4544
rect 1948 4556 1956 4564
rect 1964 4556 1972 4564
rect 2156 4556 2164 4564
rect 2236 4556 2244 4564
rect 2492 4556 2500 4564
rect 2620 4556 2628 4564
rect 2684 4556 2692 4564
rect 2908 4556 2916 4564
rect 1852 4536 1860 4544
rect 1932 4536 1940 4544
rect 2124 4536 2132 4544
rect 2172 4536 2180 4544
rect 2268 4536 2276 4544
rect 1324 4516 1332 4524
rect 1468 4516 1476 4524
rect 1660 4516 1668 4524
rect 1724 4516 1732 4524
rect 172 4496 180 4504
rect 220 4496 228 4504
rect 268 4496 276 4504
rect 444 4496 452 4504
rect 460 4496 468 4504
rect 572 4496 580 4504
rect 652 4496 660 4504
rect 716 4496 724 4504
rect 1052 4496 1060 4504
rect 1420 4496 1428 4504
rect 1500 4496 1508 4504
rect 1836 4496 1844 4504
rect 1868 4496 1876 4504
rect 1916 4516 1924 4524
rect 1996 4516 2004 4524
rect 2028 4516 2036 4524
rect 2076 4516 2084 4524
rect 2108 4516 2116 4524
rect 2188 4516 2196 4524
rect 2268 4516 2276 4524
rect 2284 4516 2292 4524
rect 2396 4516 2404 4524
rect 2428 4536 2436 4544
rect 2524 4536 2532 4544
rect 2652 4536 2660 4544
rect 2716 4536 2724 4544
rect 2732 4536 2740 4544
rect 2780 4536 2788 4544
rect 2876 4536 2884 4544
rect 3196 4556 3204 4564
rect 3756 4556 3764 4564
rect 3868 4556 3876 4564
rect 4012 4556 4020 4564
rect 4028 4556 4036 4564
rect 4092 4556 4100 4564
rect 4412 4556 4420 4564
rect 5020 4556 5028 4564
rect 5116 4556 5124 4564
rect 5452 4556 5460 4564
rect 2956 4536 2964 4544
rect 3052 4536 3060 4544
rect 3148 4536 3156 4544
rect 3228 4536 3236 4544
rect 3324 4536 3332 4544
rect 3468 4536 3476 4544
rect 3580 4536 3588 4544
rect 3740 4536 3748 4544
rect 3820 4536 3828 4544
rect 3884 4536 3892 4544
rect 3980 4536 3988 4544
rect 4028 4536 4036 4544
rect 4092 4536 4100 4544
rect 4124 4536 4132 4544
rect 4284 4536 4292 4544
rect 4316 4536 4324 4544
rect 4348 4536 4356 4544
rect 4396 4536 4404 4544
rect 4476 4536 4484 4544
rect 4540 4536 4548 4544
rect 4556 4536 4564 4544
rect 4700 4536 4708 4544
rect 4716 4536 4724 4544
rect 4828 4536 4836 4544
rect 4860 4536 4868 4544
rect 4908 4536 4916 4544
rect 5004 4536 5012 4544
rect 5084 4536 5092 4544
rect 5132 4536 5140 4544
rect 5228 4536 5236 4544
rect 5244 4536 5252 4544
rect 5276 4536 5284 4544
rect 2444 4516 2452 4524
rect 2540 4516 2548 4524
rect 2572 4516 2580 4524
rect 2668 4516 2676 4524
rect 2732 4516 2740 4524
rect 2812 4516 2820 4524
rect 2860 4516 2868 4524
rect 2940 4516 2948 4524
rect 2972 4516 2980 4524
rect 3004 4516 3012 4524
rect 3052 4516 3060 4524
rect 3244 4516 3252 4524
rect 3276 4516 3284 4524
rect 3388 4516 3396 4524
rect 3500 4516 3508 4524
rect 3612 4516 3620 4524
rect 3724 4516 3732 4524
rect 3900 4516 3908 4524
rect 3996 4516 4004 4524
rect 4140 4516 4148 4524
rect 4172 4516 4180 4524
rect 4236 4516 4244 4524
rect 5308 4532 5316 4540
rect 5404 4536 5412 4544
rect 5676 4556 5684 4564
rect 5836 4556 5844 4564
rect 6076 4556 6084 4564
rect 5564 4536 5572 4544
rect 5740 4536 5748 4544
rect 5756 4536 5764 4544
rect 5804 4536 5812 4544
rect 5820 4536 5828 4544
rect 5884 4536 5892 4544
rect 5916 4536 5924 4544
rect 5964 4536 5972 4544
rect 5980 4536 5988 4544
rect 4412 4516 4420 4524
rect 4492 4516 4500 4524
rect 4572 4516 4580 4524
rect 4716 4516 4724 4524
rect 4796 4516 4804 4524
rect 1980 4496 1988 4504
rect 2092 4496 2100 4504
rect 2220 4496 2228 4504
rect 2348 4496 2356 4504
rect 2444 4496 2452 4504
rect 2476 4496 2484 4504
rect 2556 4496 2564 4504
rect 2780 4496 2788 4504
rect 2796 4496 2804 4504
rect 2988 4496 2996 4504
rect 3084 4496 3092 4504
rect 3164 4496 3172 4504
rect 3180 4496 3188 4504
rect 3260 4496 3268 4504
rect 3356 4496 3364 4504
rect 3420 4496 3428 4504
rect 3436 4496 3444 4504
rect 3484 4496 3492 4504
rect 3548 4496 3556 4504
rect 3596 4496 3604 4504
rect 3932 4496 3940 4504
rect 3948 4496 3956 4504
rect 4076 4496 4084 4504
rect 4156 4496 4164 4504
rect 4220 4496 4228 4504
rect 4284 4496 4292 4504
rect 4508 4496 4516 4504
rect 4620 4496 4628 4504
rect 4748 4496 4756 4504
rect 4764 4496 4772 4504
rect 5372 4516 5380 4524
rect 5420 4516 5428 4524
rect 5516 4516 5524 4524
rect 5996 4532 6004 4540
rect 6076 4536 6084 4544
rect 6172 4536 6180 4544
rect 6204 4536 6212 4544
rect 5724 4516 5732 4524
rect 5788 4516 5796 4524
rect 5868 4516 5876 4524
rect 6092 4516 6100 4524
rect 4876 4496 4884 4504
rect 4972 4496 4980 4504
rect 5052 4496 5060 4504
rect 5276 4496 5284 4504
rect 5356 4496 5364 4504
rect 5596 4496 5604 4504
rect 5788 4496 5796 4504
rect 5884 4496 5892 4504
rect 5932 4496 5940 4504
rect 6172 4496 6180 4504
rect 492 4476 500 4484
rect 540 4476 548 4484
rect 940 4476 948 4484
rect 1084 4476 1092 4484
rect 1804 4476 1812 4484
rect 1980 4476 1988 4484
rect 2060 4476 2068 4484
rect 2588 4476 2596 4484
rect 2828 4476 2836 4484
rect 3020 4476 3028 4484
rect 3292 4476 3300 4484
rect 3340 4476 3348 4484
rect 3388 4476 3396 4484
rect 476 4456 484 4464
rect 556 4456 564 4464
rect 2076 4456 2084 4464
rect 2492 4456 2500 4464
rect 2812 4456 2820 4464
rect 3420 4476 3428 4484
rect 3516 4476 3524 4484
rect 3628 4476 3636 4484
rect 4188 4476 4196 4484
rect 4252 4476 4260 4484
rect 3500 4456 3508 4464
rect 684 4436 692 4444
rect 2396 4436 2404 4444
rect 2572 4436 2580 4444
rect 3068 4436 3076 4444
rect 3196 4436 3204 4444
rect 3276 4436 3284 4444
rect 6188 4436 6196 4444
rect 1566 4406 1574 4414
rect 1580 4406 1588 4414
rect 1594 4406 1602 4414
rect 4638 4406 4646 4414
rect 4652 4406 4660 4414
rect 4666 4406 4674 4414
rect 220 4376 228 4384
rect 636 4376 644 4384
rect 700 4376 708 4384
rect 844 4376 852 4384
rect 1004 4376 1012 4384
rect 1228 4376 1236 4384
rect 1308 4376 1316 4384
rect 1404 4376 1412 4384
rect 1660 4376 1668 4384
rect 1820 4376 1828 4384
rect 1900 4376 1908 4384
rect 2652 4376 2660 4384
rect 2716 4376 2724 4384
rect 2748 4376 2756 4384
rect 3052 4376 3060 4384
rect 3228 4376 3236 4384
rect 3308 4376 3316 4384
rect 3404 4376 3412 4384
rect 3564 4376 3572 4384
rect 3644 4376 3652 4384
rect 3804 4376 3812 4384
rect 3868 4376 3876 4384
rect 3948 4376 3956 4384
rect 4060 4376 4068 4384
rect 4124 4376 4132 4384
rect 4156 4376 4164 4384
rect 4188 4376 4196 4384
rect 4524 4376 4532 4384
rect 4700 4376 4708 4384
rect 4764 4376 4772 4384
rect 5100 4376 5108 4384
rect 5292 4376 5300 4384
rect 5388 4376 5396 4384
rect 5436 4376 5444 4384
rect 5500 4376 5508 4384
rect 5868 4376 5876 4384
rect 428 4356 436 4364
rect 572 4356 580 4364
rect 3164 4356 3172 4364
rect 204 4336 212 4344
rect 380 4336 388 4344
rect 444 4336 452 4344
rect 684 4336 692 4344
rect 828 4336 836 4344
rect 1148 4336 1156 4344
rect 1212 4336 1220 4344
rect 1340 4336 1348 4344
rect 1388 4336 1396 4344
rect 1676 4336 1684 4344
rect 1724 4336 1732 4344
rect 1948 4336 1956 4344
rect 2076 4336 2084 4344
rect 2396 4336 2404 4344
rect 2508 4336 2516 4344
rect 2636 4336 2644 4344
rect 2668 4336 2676 4344
rect 2972 4336 2980 4344
rect 2988 4336 2996 4344
rect 3036 4336 3044 4344
rect 3148 4336 3156 4344
rect 3212 4336 3220 4344
rect 3292 4336 3300 4344
rect 3340 4336 3348 4344
rect 3388 4336 3396 4344
rect 3548 4336 3556 4344
rect 3788 4336 3796 4344
rect 3820 4336 3828 4344
rect 3996 4336 4004 4344
rect 4044 4336 4052 4344
rect 4108 4336 4116 4344
rect 4204 4336 4212 4344
rect 5052 4336 5060 4344
rect 5084 4336 5092 4344
rect 5996 4336 6004 4344
rect 44 4316 52 4324
rect 172 4316 180 4324
rect 220 4316 228 4324
rect 316 4316 324 4324
rect 444 4316 452 4324
rect 588 4316 596 4324
rect 604 4316 612 4324
rect 716 4316 724 4324
rect 796 4316 804 4324
rect 1036 4316 1044 4324
rect 1052 4316 1060 4324
rect 1180 4316 1188 4324
rect 1244 4316 1252 4324
rect 1356 4316 1364 4324
rect 1420 4316 1428 4324
rect 1436 4316 1444 4324
rect 1516 4316 1524 4324
rect 1564 4316 1572 4324
rect 1580 4316 1588 4324
rect 1644 4316 1652 4324
rect 1692 4316 1700 4324
rect 1708 4316 1716 4324
rect 1804 4316 1812 4324
rect 1868 4316 1876 4324
rect 1980 4316 1988 4324
rect 2108 4316 2116 4324
rect 60 4296 68 4304
rect 140 4296 148 4304
rect 156 4296 164 4304
rect 220 4296 228 4304
rect 428 4296 436 4304
rect 460 4296 468 4304
rect 636 4296 644 4304
rect 700 4296 708 4304
rect 732 4296 740 4304
rect 812 4296 820 4304
rect 1004 4296 1012 4304
rect 1132 4296 1140 4304
rect 1164 4296 1172 4304
rect 1228 4296 1236 4304
rect 1260 4296 1268 4304
rect 1404 4296 1412 4304
rect 1452 4296 1460 4304
rect 1500 4296 1508 4304
rect 1660 4296 1668 4304
rect 1740 4296 1748 4304
rect 1788 4296 1796 4304
rect 1964 4296 1972 4304
rect 1996 4296 2004 4304
rect 2092 4296 2100 4304
rect 2188 4296 2196 4304
rect 2268 4296 2276 4304
rect 2364 4316 2372 4324
rect 2428 4316 2436 4324
rect 2604 4316 2612 4324
rect 2780 4316 2788 4324
rect 2956 4316 2964 4324
rect 3004 4316 3012 4324
rect 3084 4316 3092 4324
rect 3180 4316 3188 4324
rect 3244 4316 3252 4324
rect 3276 4316 3284 4324
rect 3356 4316 3364 4324
rect 3420 4316 3428 4324
rect 3500 4316 3508 4324
rect 3580 4316 3588 4324
rect 3708 4316 3716 4324
rect 3820 4316 3828 4324
rect 3916 4316 3924 4324
rect 3964 4316 3972 4324
rect 4012 4316 4020 4324
rect 4076 4316 4084 4324
rect 4252 4316 4260 4324
rect 4284 4316 4292 4324
rect 12 4276 20 4284
rect 44 4276 52 4284
rect 92 4276 100 4284
rect 316 4276 324 4284
rect 348 4276 356 4284
rect 476 4276 484 4284
rect 508 4276 516 4284
rect 556 4276 564 4284
rect 652 4276 660 4284
rect 748 4276 756 4284
rect 780 4276 788 4284
rect 908 4276 916 4284
rect 956 4276 964 4284
rect 108 4256 116 4264
rect 300 4256 308 4264
rect 364 4256 372 4264
rect 540 4256 548 4264
rect 780 4256 788 4264
rect 940 4256 948 4264
rect 1276 4276 1284 4284
rect 1324 4276 1332 4284
rect 1548 4276 1556 4284
rect 1740 4276 1748 4284
rect 1756 4276 1764 4284
rect 1852 4280 1860 4288
rect 2332 4296 2340 4304
rect 2348 4296 2356 4304
rect 2412 4296 2420 4304
rect 2444 4296 2452 4304
rect 2540 4296 2548 4304
rect 2620 4296 2628 4304
rect 2748 4296 2756 4304
rect 2892 4296 2900 4304
rect 2972 4296 2980 4304
rect 3052 4296 3060 4304
rect 3164 4296 3172 4304
rect 3228 4296 3236 4304
rect 3276 4296 3284 4304
rect 3404 4296 3412 4304
rect 3436 4296 3444 4304
rect 3484 4296 3492 4304
rect 3564 4296 3572 4304
rect 3676 4296 3684 4304
rect 3772 4296 3780 4304
rect 3836 4296 3844 4304
rect 3932 4296 3940 4304
rect 4060 4296 4068 4304
rect 4124 4296 4132 4304
rect 4220 4296 4228 4304
rect 4380 4316 4388 4324
rect 4444 4316 4452 4324
rect 4716 4316 4724 4324
rect 4844 4316 4852 4324
rect 4876 4316 4884 4324
rect 4956 4316 4964 4324
rect 5116 4316 5124 4324
rect 5244 4316 5252 4324
rect 5596 4316 5604 4324
rect 5724 4316 5732 4324
rect 5948 4316 5956 4324
rect 6060 4316 6068 4324
rect 4364 4296 4372 4304
rect 5020 4296 5028 4304
rect 5100 4296 5108 4304
rect 5500 4296 5508 4304
rect 5612 4296 5620 4304
rect 5676 4296 5684 4304
rect 5884 4296 5892 4304
rect 5996 4296 6004 4304
rect 6012 4296 6020 4304
rect 6092 4296 6100 4304
rect 6140 4296 6148 4304
rect 1868 4276 1876 4284
rect 1916 4276 1924 4284
rect 1964 4276 1972 4284
rect 2012 4276 2020 4284
rect 2204 4276 2212 4284
rect 2252 4276 2260 4284
rect 2316 4276 2324 4284
rect 2396 4276 2404 4284
rect 2460 4276 2468 4284
rect 1100 4256 1108 4264
rect 1308 4256 1316 4264
rect 1484 4256 1492 4264
rect 1532 4256 1540 4264
rect 2044 4256 2052 4264
rect 2220 4256 2228 4264
rect 2300 4256 2308 4264
rect 2556 4276 2564 4284
rect 2732 4276 2740 4284
rect 2876 4276 2884 4284
rect 3324 4276 3332 4284
rect 3452 4276 3460 4284
rect 3612 4276 3620 4284
rect 3724 4276 3732 4284
rect 3884 4276 3892 4284
rect 3932 4276 3940 4284
rect 3964 4276 3972 4284
rect 4252 4276 4260 4284
rect 4300 4276 4308 4284
rect 4428 4276 4436 4284
rect 4476 4276 4484 4284
rect 4492 4276 4500 4284
rect 4588 4276 4596 4284
rect 4732 4276 4740 4284
rect 4876 4276 4884 4284
rect 4924 4276 4932 4284
rect 4988 4276 4996 4284
rect 5004 4276 5012 4284
rect 5132 4276 5140 4284
rect 5228 4276 5236 4284
rect 5276 4276 5284 4284
rect 5324 4276 5332 4284
rect 5420 4276 5428 4284
rect 5516 4276 5524 4284
rect 5612 4276 5620 4284
rect 5628 4276 5636 4284
rect 5660 4276 5668 4284
rect 5836 4276 5844 4284
rect 5932 4276 5940 4284
rect 6108 4276 6116 4284
rect 6156 4276 6164 4284
rect 6252 4276 6260 4284
rect 2508 4256 2516 4264
rect 2588 4256 2596 4264
rect 2684 4256 2692 4264
rect 2700 4256 2708 4264
rect 2908 4256 2916 4264
rect 2924 4256 2932 4264
rect 3516 4256 3524 4264
rect 3644 4256 3652 4264
rect 3724 4256 3732 4264
rect 4172 4256 4180 4264
rect 4460 4256 4468 4264
rect 4604 4256 4612 4264
rect 4844 4256 4852 4264
rect 4940 4256 4948 4264
rect 5308 4256 5316 4264
rect 5452 4256 5460 4264
rect 5548 4256 5556 4264
rect 5852 4256 5860 4264
rect 5916 4256 5924 4264
rect 5948 4256 5956 4264
rect 6044 4256 6052 4264
rect 332 4236 340 4244
rect 492 4236 500 4244
rect 1068 4236 1076 4244
rect 1116 4236 1124 4244
rect 2028 4236 2036 4244
rect 2092 4236 2100 4244
rect 2204 4236 2212 4244
rect 2476 4236 2484 4244
rect 2572 4236 2580 4244
rect 2636 4236 2644 4244
rect 2876 4236 2884 4244
rect 2940 4236 2948 4244
rect 3628 4236 3636 4244
rect 4956 4236 4964 4244
rect 5164 4236 5172 4244
rect 5244 4236 5252 4244
rect 5644 4236 5652 4244
rect 5724 4236 5732 4244
rect 5772 4236 5780 4244
rect 5900 4236 5908 4244
rect 6060 4236 6068 4244
rect 6188 4236 6196 4244
rect 3118 4206 3126 4214
rect 3132 4206 3140 4214
rect 3146 4206 3154 4214
rect 76 4176 84 4184
rect 188 4176 196 4184
rect 252 4176 260 4184
rect 284 4176 292 4184
rect 380 4176 388 4184
rect 460 4176 468 4184
rect 588 4176 596 4184
rect 684 4176 692 4184
rect 748 4176 756 4184
rect 812 4176 820 4184
rect 1004 4176 1012 4184
rect 1020 4176 1028 4184
rect 1148 4176 1156 4184
rect 1500 4176 1508 4184
rect 1644 4176 1652 4184
rect 1740 4176 1748 4184
rect 1996 4176 2004 4184
rect 2380 4176 2388 4184
rect 2556 4176 2564 4184
rect 2700 4176 2708 4184
rect 2812 4176 2820 4184
rect 2892 4176 2900 4184
rect 3308 4176 3316 4184
rect 3388 4176 3396 4184
rect 3500 4176 3508 4184
rect 3532 4176 3540 4184
rect 3596 4176 3604 4184
rect 3692 4176 3700 4184
rect 3740 4176 3748 4184
rect 3804 4176 3812 4184
rect 3836 4176 3844 4184
rect 3916 4176 3924 4184
rect 4028 4176 4036 4184
rect 4140 4176 4148 4184
rect 4188 4176 4196 4184
rect 4252 4176 4260 4184
rect 4428 4176 4436 4184
rect 4492 4176 4500 4184
rect 4556 4176 4564 4184
rect 4684 4176 4692 4184
rect 4844 4176 4852 4184
rect 4860 4176 4868 4184
rect 5228 4176 5236 4184
rect 5292 4176 5300 4184
rect 5404 4176 5412 4184
rect 5564 4176 5572 4184
rect 5628 4176 5636 4184
rect 5836 4176 5844 4184
rect 5964 4176 5972 4184
rect 604 4156 612 4164
rect 796 4156 804 4164
rect 924 4156 932 4164
rect 940 4156 948 4164
rect 1356 4156 1364 4164
rect 1404 4156 1412 4164
rect 1580 4156 1588 4164
rect 1884 4156 1892 4164
rect 1916 4156 1924 4164
rect 2108 4156 2116 4164
rect 2124 4156 2132 4164
rect 2396 4156 2404 4164
rect 2572 4156 2580 4164
rect 3276 4156 3284 4164
rect 3548 4156 3556 4164
rect 4060 4156 4068 4164
rect 4236 4156 4244 4164
rect 4364 4156 4372 4164
rect 4476 4156 4484 4164
rect 4700 4156 4708 4164
rect 5036 4156 5044 4164
rect 5148 4156 5156 4164
rect 5532 4156 5540 4164
rect 12 4136 20 4144
rect 108 4136 116 4144
rect 124 4136 132 4144
rect 220 4136 228 4144
rect 268 4136 276 4144
rect 332 4136 340 4144
rect 348 4136 356 4144
rect 396 4136 404 4144
rect 492 4136 500 4144
rect 588 4136 596 4144
rect 636 4136 644 4144
rect 732 4136 740 4144
rect 780 4136 788 4144
rect 844 4136 852 4144
rect 860 4136 868 4144
rect 956 4136 964 4144
rect 1084 4136 1092 4144
rect 1100 4136 1108 4144
rect 1164 4136 1172 4144
rect 1212 4136 1220 4144
rect 1276 4136 1284 4144
rect 1356 4136 1364 4144
rect 1372 4136 1380 4144
rect 1420 4136 1428 4144
rect 1564 4136 1572 4144
rect 1692 4136 1700 4144
rect 1708 4136 1716 4144
rect 1804 4136 1812 4144
rect 1820 4136 1828 4144
rect 1948 4136 1956 4144
rect 2044 4136 2052 4144
rect 2060 4136 2068 4144
rect 2156 4136 2164 4144
rect 2204 4136 2212 4144
rect 2284 4136 2292 4144
rect 2364 4136 2372 4144
rect 2412 4136 2420 4144
rect 2444 4136 2452 4144
rect 2556 4136 2564 4144
rect 2652 4136 2660 4144
rect 2732 4136 2740 4144
rect 2860 4136 2868 4144
rect 2940 4136 2948 4144
rect 3180 4136 3188 4144
rect 3228 4136 3236 4144
rect 3244 4136 3252 4144
rect 3420 4136 3428 4144
rect 3436 4136 3444 4144
rect 3564 4136 3572 4144
rect 3612 4136 3620 4144
rect 3644 4136 3652 4144
rect 3708 4136 3716 4144
rect 3756 4136 3764 4144
rect 3820 4136 3828 4144
rect 3868 4136 3876 4144
rect 332 4116 340 4124
rect 588 4116 596 4124
rect 732 4116 740 4124
rect 876 4116 884 4124
rect 972 4116 980 4124
rect 1116 4116 1124 4124
rect 1228 4116 1236 4124
rect 1244 4116 1252 4124
rect 1292 4116 1300 4124
rect 1324 4116 1332 4124
rect 1436 4116 1444 4124
rect 1676 4116 1684 4124
rect 1836 4116 1844 4124
rect 1916 4116 1924 4124
rect 2076 4116 2084 4124
rect 2156 4116 2164 4124
rect 2204 4116 2212 4124
rect 2236 4116 2244 4124
rect 2300 4116 2308 4124
rect 2428 4116 2436 4124
rect 2540 4116 2548 4124
rect 2684 4116 2692 4124
rect 2748 4116 2756 4124
rect 2780 4116 2788 4124
rect 2812 4116 2820 4124
rect 2940 4116 2948 4124
rect 2972 4116 2980 4124
rect 3020 4116 3028 4124
rect 3084 4116 3092 4124
rect 3212 4116 3220 4124
rect 3324 4116 3332 4124
rect 3388 4116 3396 4124
rect 236 4096 244 4104
rect 284 4096 292 4104
rect 380 4096 388 4104
rect 684 4096 692 4104
rect 700 4096 708 4104
rect 812 4096 820 4104
rect 908 4096 916 4104
rect 1052 4096 1060 4104
rect 1196 4096 1204 4104
rect 1260 4096 1268 4104
rect 1324 4096 1332 4104
rect 1404 4096 1412 4104
rect 1468 4096 1476 4104
rect 1644 4096 1652 4104
rect 1868 4096 1876 4104
rect 1996 4096 2004 4104
rect 2108 4096 2116 4104
rect 2220 4096 2228 4104
rect 2332 4096 2340 4104
rect 2460 4096 2468 4104
rect 2652 4096 2660 4104
rect 2684 4096 2692 4104
rect 2780 4096 2788 4104
rect 2796 4096 2804 4104
rect 2892 4096 2900 4104
rect 2956 4096 2964 4104
rect 3004 4096 3012 4104
rect 3068 4096 3076 4104
rect 3340 4096 3348 4104
rect 3404 4096 3412 4104
rect 3468 4096 3476 4104
rect 3516 4116 3524 4124
rect 3564 4116 3572 4124
rect 3628 4116 3636 4124
rect 3660 4116 3668 4124
rect 3772 4116 3780 4124
rect 3932 4116 3940 4124
rect 3980 4136 3988 4144
rect 4172 4136 4180 4144
rect 4220 4136 4228 4144
rect 4284 4136 4292 4144
rect 4380 4136 4388 4144
rect 4396 4136 4404 4144
rect 4460 4136 4468 4144
rect 4524 4136 4532 4144
rect 4572 4136 4580 4144
rect 4780 4136 4788 4144
rect 4908 4136 4916 4144
rect 5004 4136 5012 4144
rect 5116 4136 5124 4144
rect 5164 4136 5172 4144
rect 5180 4136 5188 4144
rect 5244 4136 5252 4144
rect 5308 4136 5316 4144
rect 5356 4136 5364 4144
rect 5756 4156 5764 4164
rect 5724 4136 5732 4144
rect 6044 4136 6052 4144
rect 6156 4136 6164 4144
rect 6172 4136 6180 4144
rect 3996 4116 4004 4124
rect 4108 4116 4116 4124
rect 4332 4116 4340 4124
rect 4412 4116 4420 4124
rect 4604 4116 4612 4124
rect 4780 4116 4788 4124
rect 4892 4116 4900 4124
rect 4956 4116 4964 4124
rect 4988 4116 4996 4124
rect 5052 4116 5060 4124
rect 5100 4116 5108 4124
rect 5164 4116 5172 4124
rect 5196 4116 5204 4124
rect 5244 4116 5252 4124
rect 5324 4116 5332 4124
rect 5404 4116 5412 4124
rect 5452 4116 5460 4124
rect 5500 4116 5508 4124
rect 5596 4116 5604 4124
rect 5676 4116 5684 4124
rect 5708 4116 5716 4124
rect 5756 4116 5764 4124
rect 5820 4116 5828 4124
rect 5884 4116 5892 4124
rect 5964 4116 5972 4124
rect 6028 4116 6036 4124
rect 6108 4116 6116 4124
rect 6172 4116 6180 4124
rect 3708 4096 3716 4104
rect 3740 4096 3748 4104
rect 3804 4096 3812 4104
rect 3852 4096 3860 4104
rect 4124 4096 4132 4104
rect 4140 4096 4148 4104
rect 4252 4096 4260 4104
rect 4348 4096 4356 4104
rect 4492 4096 4500 4104
rect 4540 4096 4548 4104
rect 4588 4096 4596 4104
rect 4764 4096 4772 4104
rect 4844 4096 4852 4104
rect 4860 4096 4868 4104
rect 4972 4096 4980 4104
rect 5052 4096 5060 4104
rect 5292 4096 5300 4104
rect 5356 4096 5364 4104
rect 5420 4096 5428 4104
rect 5692 4096 5700 4104
rect 5804 4096 5812 4104
rect 5868 4096 5876 4104
rect 5996 4096 6004 4104
rect 6108 4096 6116 4104
rect 6124 4096 6132 4104
rect 6220 4096 6228 4104
rect 1516 4076 1524 4084
rect 1980 4076 1988 4084
rect 2252 4076 2260 4084
rect 2700 4076 2708 4084
rect 2828 4076 2836 4084
rect 2988 4076 2996 4084
rect 3100 4076 3108 4084
rect 3276 4076 3284 4084
rect 3308 4076 3316 4084
rect 3372 4076 3380 4084
rect 4092 4076 4100 4084
rect 4316 4076 4324 4084
rect 4620 4076 4628 4084
rect 4668 4076 4676 4084
rect 4940 4076 4948 4084
rect 5388 4076 5396 4084
rect 5404 4076 5412 4084
rect 5660 4076 5668 4084
rect 5884 4076 5892 4084
rect 5900 4076 5908 4084
rect 5948 4076 5956 4084
rect 2236 4056 2244 4064
rect 3052 4056 3060 4064
rect 4108 4056 4116 4064
rect 4956 4056 4964 4064
rect 5484 4056 5492 4064
rect 828 4036 836 4044
rect 1836 4036 1844 4044
rect 1900 4036 1908 4044
rect 2716 4036 2724 4044
rect 2748 4036 2756 4044
rect 3164 4036 3172 4044
rect 4044 4036 4052 4044
rect 4332 4036 4340 4044
rect 5676 4036 5684 4044
rect 5884 4036 5892 4044
rect 5964 4036 5972 4044
rect 6028 4036 6036 4044
rect 6076 4036 6084 4044
rect 6188 4036 6196 4044
rect 1566 4006 1574 4014
rect 1580 4006 1588 4014
rect 1594 4006 1602 4014
rect 4638 4006 4646 4014
rect 4652 4006 4660 4014
rect 4666 4006 4674 4014
rect 76 3976 84 3984
rect 188 3976 196 3984
rect 444 3976 452 3984
rect 572 3976 580 3984
rect 716 3976 724 3984
rect 796 3976 804 3984
rect 844 3976 852 3984
rect 908 3976 916 3984
rect 1100 3976 1108 3984
rect 1196 3976 1204 3984
rect 1324 3976 1332 3984
rect 1500 3976 1508 3984
rect 1692 3976 1700 3984
rect 1964 3976 1972 3984
rect 1996 3976 2004 3984
rect 2220 3976 2228 3984
rect 2236 3976 2244 3984
rect 2652 3976 2660 3984
rect 2684 3976 2692 3984
rect 2812 3976 2820 3984
rect 2924 3976 2932 3984
rect 2972 3976 2980 3984
rect 3132 3976 3140 3984
rect 3244 3976 3252 3984
rect 3276 3976 3284 3984
rect 3340 3976 3348 3984
rect 3692 3976 3700 3984
rect 3740 3976 3748 3984
rect 4140 3976 4148 3984
rect 4204 3976 4212 3984
rect 4316 3976 4324 3984
rect 4396 3976 4404 3984
rect 4444 3976 4452 3984
rect 4476 3976 4484 3984
rect 4556 3976 4564 3984
rect 4780 3976 4788 3984
rect 4908 3976 4916 3984
rect 5004 3976 5012 3984
rect 5036 3976 5044 3984
rect 5132 3976 5140 3984
rect 5468 3976 5476 3984
rect 5612 3976 5620 3984
rect 6124 3976 6132 3984
rect 6140 3976 6148 3984
rect 1036 3956 1044 3964
rect 1436 3956 1444 3964
rect 1916 3956 1924 3964
rect 3420 3956 3428 3964
rect 3484 3956 3492 3964
rect 4060 3956 4068 3964
rect 204 3936 212 3944
rect 364 3936 372 3944
rect 556 3936 564 3944
rect 700 3936 708 3944
rect 732 3936 740 3944
rect 972 3936 980 3944
rect 1148 3936 1156 3944
rect 2204 3936 2212 3944
rect 2332 3936 2340 3944
rect 2764 3936 2772 3944
rect 2796 3936 2804 3944
rect 2844 3936 2852 3944
rect 2956 3936 2964 3944
rect 3404 3936 3412 3944
rect 3468 3936 3476 3944
rect 3676 3936 3684 3944
rect 3724 3936 3732 3944
rect 3916 3936 3924 3944
rect 3980 3936 3988 3944
rect 4044 3936 4052 3944
rect 4188 3936 4196 3944
rect 4252 3936 4260 3944
rect 4300 3936 4308 3944
rect 4428 3936 4436 3944
rect 4860 3936 4868 3944
rect 4892 3936 4900 3944
rect 4988 3936 4996 3944
rect 5740 3936 5748 3944
rect 5804 3936 5812 3944
rect 5868 3936 5876 3944
rect 5884 3936 5892 3944
rect 5980 3936 5988 3944
rect 6028 3936 6036 3944
rect 6060 3936 6068 3944
rect 124 3916 132 3924
rect 236 3916 244 3924
rect 268 3916 276 3924
rect 508 3916 516 3924
rect 620 3916 628 3924
rect 668 3916 676 3924
rect 876 3916 884 3924
rect 940 3916 948 3924
rect 1052 3916 1060 3924
rect 1068 3916 1076 3924
rect 1164 3916 1172 3924
rect 140 3896 148 3904
rect 156 3896 164 3904
rect 204 3896 212 3904
rect 252 3896 260 3904
rect 364 3896 372 3904
rect 396 3896 404 3904
rect 412 3896 420 3904
rect 476 3896 484 3904
rect 540 3896 548 3904
rect 652 3896 660 3904
rect 700 3896 708 3904
rect 796 3896 804 3904
rect 908 3896 916 3904
rect 956 3896 964 3904
rect 972 3896 980 3904
rect 1100 3896 1108 3904
rect 1196 3896 1204 3904
rect 1244 3916 1252 3924
rect 1420 3916 1428 3924
rect 2156 3916 2164 3924
rect 2172 3916 2180 3924
rect 2300 3916 2308 3924
rect 2604 3916 2612 3924
rect 2620 3916 2628 3924
rect 2748 3916 2756 3924
rect 2764 3916 2772 3924
rect 1276 3896 1284 3904
rect 1324 3896 1332 3904
rect 1612 3896 1620 3904
rect 1660 3896 1668 3904
rect 1820 3896 1828 3904
rect 1964 3896 1972 3904
rect 2044 3896 2052 3904
rect 2156 3896 2164 3904
rect 2188 3896 2196 3904
rect 2284 3896 2292 3904
rect 2540 3896 2548 3904
rect 2652 3896 2660 3904
rect 2780 3896 2788 3904
rect 3004 3916 3012 3924
rect 3036 3916 3044 3924
rect 3068 3916 3076 3924
rect 3148 3916 3156 3924
rect 3308 3916 3316 3924
rect 3372 3916 3380 3924
rect 3436 3916 3444 3924
rect 3500 3916 3508 3924
rect 3516 3916 3524 3924
rect 3548 3916 3556 3924
rect 3644 3916 3652 3924
rect 3756 3916 3764 3924
rect 3884 3916 3892 3924
rect 3948 3916 3956 3924
rect 4012 3916 4020 3924
rect 4076 3916 4084 3924
rect 4092 3916 4100 3924
rect 4156 3916 4164 3924
rect 4220 3916 4228 3924
rect 4332 3916 4340 3924
rect 4460 3916 4468 3924
rect 2876 3896 2884 3904
rect 2972 3896 2980 3904
rect 3052 3896 3060 3904
rect 3100 3896 3108 3904
rect 3196 3896 3204 3904
rect 3244 3896 3252 3904
rect 3276 3896 3284 3904
rect 3340 3896 3348 3904
rect 3420 3896 3428 3904
rect 3484 3896 3492 3904
rect 3548 3896 3556 3904
rect 3580 3896 3588 3904
rect 3628 3896 3636 3904
rect 3660 3896 3668 3904
rect 3740 3896 3748 3904
rect 3772 3896 3780 3904
rect 3852 3896 3860 3904
rect 3900 3896 3908 3904
rect 3916 3896 3924 3904
rect 3996 3896 4004 3904
rect 4060 3896 4068 3904
rect 4108 3896 4116 3904
rect 4172 3896 4180 3904
rect 4236 3896 4244 3904
rect 4268 3896 4276 3904
rect 4316 3896 4324 3904
rect 4348 3896 4356 3904
rect 4444 3896 4452 3904
rect 4508 3896 4516 3904
rect 4572 3896 4580 3904
rect 4588 3896 4596 3904
rect 4828 3916 4836 3924
rect 5020 3916 5028 3924
rect 5212 3916 5220 3924
rect 5244 3916 5252 3924
rect 5324 3916 5332 3924
rect 5580 3916 5588 3924
rect 5660 3916 5668 3924
rect 5692 3916 5700 3924
rect 5708 3916 5716 3924
rect 5836 3916 5844 3924
rect 5900 3916 5908 3924
rect 6172 3916 6180 3924
rect 4908 3896 4916 3904
rect 5004 3896 5012 3904
rect 5100 3896 5108 3904
rect 5132 3896 5140 3904
rect 5164 3896 5172 3904
rect 5196 3896 5204 3904
rect 5324 3896 5332 3904
rect 5564 3896 5572 3904
rect 5612 3896 5620 3904
rect 5660 3896 5668 3904
rect 5820 3896 5828 3904
rect 5884 3896 5892 3904
rect 5964 3896 5972 3904
rect 6044 3896 6052 3904
rect 6076 3896 6084 3904
rect 6220 3896 6228 3904
rect 12 3876 20 3884
rect 108 3876 116 3884
rect 172 3876 180 3884
rect 284 3876 292 3884
rect 412 3876 420 3884
rect 588 3876 596 3884
rect 636 3876 644 3884
rect 812 3876 820 3884
rect 828 3876 836 3884
rect 892 3876 900 3884
rect 956 3876 964 3884
rect 1020 3876 1028 3884
rect 1116 3876 1124 3884
rect 1132 3876 1140 3884
rect 1292 3876 1300 3884
rect 1340 3876 1348 3884
rect 1372 3876 1380 3884
rect 1468 3876 1476 3884
rect 1516 3876 1524 3884
rect 284 3856 292 3864
rect 508 3856 516 3864
rect 636 3856 644 3864
rect 748 3856 756 3864
rect 1388 3856 1396 3864
rect 1420 3856 1428 3864
rect 1452 3856 1460 3864
rect 1708 3876 1716 3884
rect 1804 3876 1812 3884
rect 1884 3876 1892 3884
rect 2060 3876 2068 3884
rect 2268 3876 2276 3884
rect 2348 3876 2356 3884
rect 2396 3876 2404 3884
rect 2492 3876 2500 3884
rect 2556 3876 2564 3884
rect 2572 3876 2580 3884
rect 2668 3876 2676 3884
rect 2716 3876 2724 3884
rect 2828 3876 2836 3884
rect 2892 3876 2900 3884
rect 3196 3876 3204 3884
rect 3244 3876 3252 3884
rect 3324 3876 3332 3884
rect 3564 3876 3572 3884
rect 3596 3876 3604 3884
rect 3788 3876 3796 3884
rect 3836 3876 3844 3884
rect 3900 3876 3908 3884
rect 3980 3876 3988 3884
rect 4364 3876 4372 3884
rect 4524 3876 4532 3884
rect 4652 3876 4660 3884
rect 4716 3876 4724 3884
rect 4828 3876 4836 3884
rect 4860 3876 4868 3884
rect 5148 3876 5156 3884
rect 5244 3876 5252 3884
rect 5292 3876 5300 3884
rect 5356 3876 5364 3884
rect 5388 3876 5396 3884
rect 5420 3876 5428 3884
rect 5516 3876 5524 3884
rect 5628 3876 5636 3884
rect 5644 3876 5652 3884
rect 5708 3876 5716 3884
rect 5740 3876 5748 3884
rect 6076 3876 6084 3884
rect 6236 3876 6244 3884
rect 1628 3856 1636 3864
rect 1852 3856 1860 3864
rect 1868 3856 1876 3864
rect 1932 3856 1940 3864
rect 2076 3856 2084 3864
rect 2236 3856 2244 3864
rect 2380 3856 2388 3864
rect 2700 3856 2708 3864
rect 2924 3856 2932 3864
rect 3004 3856 3012 3864
rect 3212 3856 3220 3864
rect 3628 3856 3636 3864
rect 3820 3856 3828 3864
rect 4396 3856 4404 3864
rect 4492 3856 4500 3864
rect 4556 3856 4564 3864
rect 4604 3856 4612 3864
rect 4956 3856 4964 3864
rect 5052 3856 5060 3864
rect 5068 3856 5076 3864
rect 5100 3856 5108 3864
rect 5308 3856 5316 3864
rect 5372 3856 5380 3864
rect 5532 3856 5540 3864
rect 5548 3856 5556 3864
rect 5772 3856 5780 3864
rect 5932 3856 5940 3864
rect 6124 3856 6132 3864
rect 6156 3856 6164 3864
rect 1436 3836 1444 3844
rect 1772 3836 1780 3844
rect 2460 3836 2468 3844
rect 2508 3836 2516 3844
rect 2604 3836 2612 3844
rect 2748 3836 2756 3844
rect 4636 3836 4644 3844
rect 5196 3836 5204 3844
rect 5820 3836 5828 3844
rect 5884 3836 5892 3844
rect 5964 3836 5972 3844
rect 6044 3836 6052 3844
rect 6108 3836 6116 3844
rect 3118 3806 3126 3814
rect 3132 3806 3140 3814
rect 3146 3806 3154 3814
rect 44 3776 52 3784
rect 172 3776 180 3784
rect 204 3776 212 3784
rect 236 3776 244 3784
rect 380 3776 388 3784
rect 412 3776 420 3784
rect 540 3776 548 3784
rect 604 3776 612 3784
rect 668 3776 676 3784
rect 748 3776 756 3784
rect 828 3776 836 3784
rect 892 3776 900 3784
rect 1084 3776 1092 3784
rect 1148 3776 1156 3784
rect 1628 3776 1636 3784
rect 1836 3776 1844 3784
rect 1980 3776 1988 3784
rect 2172 3776 2180 3784
rect 2236 3776 2244 3784
rect 2396 3776 2404 3784
rect 2636 3776 2644 3784
rect 2716 3776 2724 3784
rect 2780 3776 2788 3784
rect 2876 3776 2884 3784
rect 2956 3776 2964 3784
rect 3244 3776 3252 3784
rect 3356 3776 3364 3784
rect 3452 3776 3460 3784
rect 3516 3776 3524 3784
rect 3580 3776 3588 3784
rect 3644 3776 3652 3784
rect 3692 3776 3700 3784
rect 3724 3776 3732 3784
rect 3820 3776 3828 3784
rect 3900 3776 3908 3784
rect 4044 3776 4052 3784
rect 4188 3776 4196 3784
rect 4284 3776 4292 3784
rect 4332 3776 4340 3784
rect 4396 3776 4404 3784
rect 4428 3776 4436 3784
rect 4460 3776 4468 3784
rect 4508 3776 4516 3784
rect 4604 3776 4612 3784
rect 4732 3776 4740 3784
rect 4908 3776 4916 3784
rect 4988 3776 4996 3784
rect 5004 3776 5012 3784
rect 5084 3776 5092 3784
rect 5132 3776 5140 3784
rect 5324 3776 5332 3784
rect 5372 3776 5380 3784
rect 5436 3776 5444 3784
rect 5500 3776 5508 3784
rect 5676 3776 5684 3784
rect 5692 3776 5700 3784
rect 5852 3776 5860 3784
rect 6124 3776 6132 3784
rect 124 3756 132 3764
rect 396 3756 404 3764
rect 652 3756 660 3764
rect 732 3756 740 3764
rect 1020 3756 1028 3764
rect 1052 3756 1060 3764
rect 12 3736 20 3744
rect 140 3736 148 3744
rect 188 3736 196 3744
rect 284 3736 292 3744
rect 300 3736 308 3744
rect 460 3736 468 3744
rect 476 3736 484 3744
rect 508 3736 516 3744
rect 556 3736 564 3744
rect 572 3736 580 3744
rect 620 3736 628 3744
rect 732 3736 740 3744
rect 780 3736 788 3744
rect 796 3732 804 3740
rect 844 3736 852 3744
rect 908 3736 916 3744
rect 956 3736 964 3744
rect 1132 3756 1140 3764
rect 1196 3756 1204 3764
rect 1852 3756 1860 3764
rect 2044 3756 2052 3764
rect 2060 3756 2068 3764
rect 2380 3756 2388 3764
rect 2508 3756 2516 3764
rect 1100 3736 1108 3744
rect 1164 3736 1172 3744
rect 1212 3736 1220 3744
rect 1308 3736 1316 3744
rect 268 3716 276 3724
rect 316 3716 324 3724
rect 332 3716 340 3724
rect 364 3716 372 3724
rect 476 3716 484 3724
rect 220 3696 228 3704
rect 348 3696 356 3704
rect 412 3696 420 3704
rect 476 3696 484 3704
rect 524 3696 532 3704
rect 604 3696 612 3704
rect 652 3696 660 3704
rect 716 3716 724 3724
rect 764 3716 772 3724
rect 844 3716 852 3724
rect 956 3716 964 3724
rect 1020 3716 1028 3724
rect 1116 3716 1124 3724
rect 1164 3716 1172 3724
rect 1356 3736 1364 3744
rect 1388 3736 1396 3744
rect 1436 3736 1444 3744
rect 1484 3736 1492 3744
rect 1548 3736 1556 3744
rect 1644 3736 1652 3744
rect 1740 3736 1748 3744
rect 1804 3736 1812 3744
rect 1868 3736 1876 3744
rect 1884 3732 1892 3740
rect 1932 3736 1940 3744
rect 1996 3736 2004 3744
rect 2092 3736 2100 3744
rect 2140 3736 2148 3744
rect 2188 3736 2196 3744
rect 2268 3736 2276 3744
rect 2412 3736 2420 3744
rect 2476 3736 2484 3744
rect 2652 3736 2660 3744
rect 2828 3756 2836 3764
rect 2940 3756 2948 3764
rect 3052 3756 3060 3764
rect 3212 3756 3220 3764
rect 2732 3736 2740 3744
rect 2764 3736 2772 3744
rect 2844 3736 2852 3744
rect 2892 3736 2900 3744
rect 2924 3736 2932 3744
rect 2972 3736 2980 3744
rect 3004 3736 3012 3744
rect 3068 3736 3076 3744
rect 3436 3756 3444 3764
rect 3596 3756 3604 3764
rect 3612 3756 3620 3764
rect 3628 3756 3636 3764
rect 3708 3756 3716 3764
rect 4476 3756 4484 3764
rect 4748 3756 4756 3764
rect 4844 3756 4852 3764
rect 5052 3756 5060 3764
rect 5612 3756 5620 3764
rect 5708 3756 5716 3764
rect 5740 3756 5748 3764
rect 5772 3756 5780 3764
rect 3260 3736 3268 3744
rect 3292 3736 3300 3744
rect 3340 3736 3348 3744
rect 3420 3736 3428 3744
rect 3468 3736 3476 3744
rect 3532 3736 3540 3744
rect 3564 3736 3572 3744
rect 3756 3736 3764 3744
rect 3772 3736 3780 3744
rect 3788 3732 3796 3740
rect 3836 3736 3844 3744
rect 3932 3736 3940 3744
rect 3948 3736 3956 3744
rect 3980 3736 3988 3744
rect 4220 3736 4228 3744
rect 4236 3736 4244 3744
rect 4300 3736 4308 3744
rect 4332 3736 4340 3744
rect 4412 3736 4420 3744
rect 4588 3736 4596 3744
rect 4812 3736 4820 3744
rect 4860 3736 4868 3744
rect 4908 3736 4916 3744
rect 4940 3736 4948 3744
rect 5084 3736 5092 3744
rect 5116 3736 5124 3744
rect 5244 3736 5252 3744
rect 5260 3736 5268 3744
rect 5356 3736 5364 3744
rect 5420 3736 5428 3744
rect 5468 3732 5476 3740
rect 5484 3736 5492 3744
rect 5548 3736 5556 3744
rect 5564 3736 5572 3744
rect 5628 3736 5636 3744
rect 5708 3736 5716 3744
rect 5868 3756 5876 3764
rect 5884 3756 5892 3764
rect 5980 3756 5988 3764
rect 6012 3756 6020 3764
rect 6108 3756 6116 3764
rect 6220 3756 6228 3764
rect 5804 3736 5812 3744
rect 6012 3736 6020 3744
rect 6108 3736 6116 3744
rect 6140 3736 6148 3744
rect 6156 3736 6164 3744
rect 6220 3736 6228 3744
rect 1340 3716 1348 3724
rect 1372 3716 1380 3724
rect 1500 3716 1508 3724
rect 1548 3716 1556 3724
rect 1772 3716 1780 3724
rect 1788 3716 1796 3724
rect 1820 3716 1828 3724
rect 1948 3716 1956 3724
rect 2012 3716 2020 3724
rect 2092 3716 2100 3724
rect 2204 3716 2212 3724
rect 2284 3716 2292 3724
rect 2348 3716 2356 3724
rect 2508 3716 2516 3724
rect 2572 3716 2580 3724
rect 2748 3716 2756 3724
rect 3020 3716 3028 3724
rect 3084 3716 3092 3724
rect 3180 3716 3188 3724
rect 3276 3716 3284 3724
rect 3484 3716 3492 3724
rect 3532 3716 3540 3724
rect 3676 3716 3684 3724
rect 3996 3716 4004 3724
rect 4012 3716 4020 3724
rect 4076 3716 4084 3724
rect 4108 3716 4116 3724
rect 4156 3716 4164 3724
rect 4252 3716 4260 3724
rect 4364 3716 4372 3724
rect 4572 3716 4580 3724
rect 4636 3716 4644 3724
rect 4716 3716 4724 3724
rect 4780 3716 4788 3724
rect 5164 3716 5172 3724
rect 5228 3716 5236 3724
rect 5404 3716 5412 3724
rect 5532 3716 5540 3724
rect 5580 3716 5588 3724
rect 5644 3716 5652 3724
rect 5756 3716 5764 3724
rect 5820 3716 5828 3724
rect 5932 3716 5940 3724
rect 6060 3716 6068 3724
rect 6156 3716 6164 3724
rect 892 3696 900 3704
rect 940 3696 948 3704
rect 1004 3696 1012 3704
rect 1372 3696 1380 3704
rect 1388 3696 1396 3704
rect 1420 3696 1428 3704
rect 1436 3696 1444 3704
rect 1468 3696 1476 3704
rect 1532 3696 1540 3704
rect 1580 3696 1588 3704
rect 1628 3696 1636 3704
rect 1756 3696 1764 3704
rect 1980 3696 1988 3704
rect 2124 3696 2132 3704
rect 2188 3696 2196 3704
rect 2300 3696 2308 3704
rect 2364 3696 2372 3704
rect 2444 3696 2452 3704
rect 2492 3696 2500 3704
rect 2556 3696 2564 3704
rect 2620 3696 2628 3704
rect 2876 3696 2884 3704
rect 2924 3696 2932 3704
rect 3004 3696 3012 3704
rect 3084 3696 3092 3704
rect 3116 3696 3124 3704
rect 3292 3696 3300 3704
rect 3388 3696 3396 3704
rect 3500 3696 3508 3704
rect 3724 3696 3732 3704
rect 3980 3696 3988 3704
rect 4044 3696 4052 3704
rect 4060 3696 4068 3704
rect 4172 3696 4180 3704
rect 4188 3696 4196 3704
rect 4332 3696 4340 3704
rect 4444 3696 4452 3704
rect 4492 3696 4500 3704
rect 4540 3696 4548 3704
rect 4892 3696 4900 3704
rect 4908 3696 4916 3704
rect 5004 3696 5012 3704
rect 5084 3696 5092 3704
rect 5196 3696 5204 3704
rect 5612 3696 5620 3704
rect 5852 3696 5860 3704
rect 5948 3696 5956 3704
rect 5964 3696 5972 3704
rect 2108 3676 2116 3684
rect 2268 3676 2276 3684
rect 2332 3676 2340 3684
rect 2492 3676 2500 3684
rect 2524 3676 2532 3684
rect 2588 3676 2596 3684
rect 3308 3676 3316 3684
rect 4092 3676 4100 3684
rect 4140 3676 4148 3684
rect 5916 3676 5924 3684
rect 6076 3676 6084 3684
rect 4076 3656 4084 3664
rect 4156 3656 4164 3664
rect 924 3636 932 3644
rect 1180 3636 1188 3644
rect 1276 3636 1284 3644
rect 1452 3636 1460 3644
rect 1708 3636 1716 3644
rect 2348 3636 2356 3644
rect 2604 3636 2612 3644
rect 3196 3636 3204 3644
rect 5932 3636 5940 3644
rect 1566 3606 1574 3614
rect 1580 3606 1588 3614
rect 1594 3606 1602 3614
rect 4638 3606 4646 3614
rect 4652 3606 4660 3614
rect 4666 3606 4674 3614
rect 76 3576 84 3584
rect 172 3576 180 3584
rect 300 3576 308 3584
rect 364 3576 372 3584
rect 412 3576 420 3584
rect 492 3576 500 3584
rect 556 3576 564 3584
rect 636 3576 644 3584
rect 700 3576 708 3584
rect 796 3576 804 3584
rect 1244 3576 1252 3584
rect 1340 3576 1348 3584
rect 1372 3576 1380 3584
rect 1660 3576 1668 3584
rect 2044 3576 2052 3584
rect 2428 3576 2436 3584
rect 2508 3576 2516 3584
rect 2652 3576 2660 3584
rect 3084 3576 3092 3584
rect 3228 3576 3236 3584
rect 3356 3576 3364 3584
rect 3436 3576 3444 3584
rect 3468 3576 3476 3584
rect 3580 3576 3588 3584
rect 3740 3576 3748 3584
rect 3836 3576 3844 3584
rect 3964 3576 3972 3584
rect 4204 3576 4212 3584
rect 4252 3576 4260 3584
rect 4396 3576 4404 3584
rect 4460 3576 4468 3584
rect 4508 3576 4516 3584
rect 4604 3576 4612 3584
rect 4956 3576 4964 3584
rect 5116 3576 5124 3584
rect 5164 3576 5172 3584
rect 5340 3576 5348 3584
rect 5436 3576 5444 3584
rect 5772 3576 5780 3584
rect 5836 3576 5844 3584
rect 5868 3576 5876 3584
rect 5996 3576 6004 3584
rect 2188 3556 2196 3564
rect 4364 3556 4372 3564
rect 4828 3556 4836 3564
rect 5516 3556 5524 3564
rect 140 3536 148 3544
rect 460 3536 468 3544
rect 940 3536 948 3544
rect 956 3536 964 3544
rect 1260 3536 1268 3544
rect 1356 3536 1364 3544
rect 1372 3536 1380 3544
rect 1612 3536 1620 3544
rect 1788 3536 1796 3544
rect 2172 3536 2180 3544
rect 2348 3536 2356 3544
rect 2796 3536 2804 3544
rect 3036 3536 3044 3544
rect 3100 3536 3108 3544
rect 3244 3536 3252 3544
rect 3692 3536 3700 3544
rect 3724 3536 3732 3544
rect 4300 3536 4308 3544
rect 4412 3536 4420 3544
rect 4476 3536 4484 3544
rect 4924 3536 4932 3544
rect 5228 3536 5236 3544
rect 5724 3536 5732 3544
rect 5820 3536 5828 3544
rect 5884 3536 5892 3544
rect 6188 3536 6196 3544
rect 172 3496 180 3504
rect 220 3516 228 3524
rect 332 3516 340 3524
rect 428 3516 436 3524
rect 764 3516 772 3524
rect 828 3516 836 3524
rect 908 3516 916 3524
rect 1148 3516 1156 3524
rect 1212 3516 1220 3524
rect 1356 3516 1364 3524
rect 1468 3516 1476 3524
rect 1644 3516 1652 3524
rect 1788 3516 1796 3524
rect 1932 3514 1940 3522
rect 2076 3516 2084 3524
rect 2140 3516 2148 3524
rect 2204 3516 2212 3524
rect 2348 3516 2356 3524
rect 2540 3516 2548 3524
rect 268 3496 276 3504
rect 332 3496 340 3504
rect 460 3496 468 3504
rect 476 3496 484 3504
rect 556 3496 564 3504
rect 588 3496 596 3504
rect 652 3496 660 3504
rect 716 3496 724 3504
rect 780 3496 788 3504
rect 796 3496 804 3504
rect 828 3496 836 3504
rect 924 3496 932 3504
rect 1036 3496 1044 3504
rect 1116 3496 1124 3504
rect 1180 3496 1188 3504
rect 1244 3496 1252 3504
rect 1292 3496 1300 3504
rect 1372 3496 1380 3504
rect 1420 3496 1428 3504
rect 1436 3496 1444 3504
rect 1484 3496 1492 3504
rect 1596 3496 1604 3504
rect 1612 3496 1620 3504
rect 1708 3496 1716 3504
rect 108 3476 116 3484
rect 156 3476 164 3484
rect 268 3476 276 3484
rect 284 3476 292 3484
rect 492 3476 500 3484
rect 540 3476 548 3484
rect 604 3476 612 3484
rect 780 3476 788 3484
rect 860 3476 868 3484
rect 876 3476 884 3484
rect 1052 3476 1060 3484
rect 1164 3476 1172 3484
rect 1308 3476 1316 3484
rect 1420 3476 1428 3484
rect 1500 3476 1508 3484
rect 1564 3476 1572 3484
rect 1692 3476 1700 3484
rect 1804 3496 1812 3504
rect 1852 3496 1860 3504
rect 1884 3496 1892 3504
rect 1964 3496 1972 3504
rect 2044 3496 2052 3504
rect 2076 3496 2084 3504
rect 2188 3496 2196 3504
rect 2220 3496 2228 3504
rect 2284 3496 2292 3504
rect 2364 3496 2372 3504
rect 2412 3496 2420 3504
rect 2444 3496 2452 3504
rect 2524 3496 2532 3504
rect 2588 3516 2596 3524
rect 2684 3516 2692 3524
rect 2764 3516 2772 3524
rect 3004 3516 3012 3524
rect 3068 3516 3076 3524
rect 3276 3516 3284 3524
rect 3292 3516 3300 3524
rect 2748 3496 2756 3504
rect 2780 3496 2788 3504
rect 2988 3496 2996 3504
rect 3020 3496 3028 3504
rect 3084 3496 3092 3504
rect 3212 3496 3220 3504
rect 3260 3496 3268 3504
rect 3292 3496 3300 3504
rect 3324 3496 3332 3504
rect 3388 3496 3396 3504
rect 3468 3496 3476 3504
rect 3596 3516 3604 3524
rect 3612 3516 3620 3524
rect 3756 3516 3764 3524
rect 4076 3516 4084 3524
rect 4156 3516 4164 3524
rect 4268 3516 4276 3524
rect 4332 3516 4340 3524
rect 4380 3516 4388 3524
rect 4444 3516 4452 3524
rect 4764 3516 4772 3524
rect 4892 3516 4900 3524
rect 5084 3516 5092 3524
rect 5196 3516 5204 3524
rect 5212 3516 5220 3524
rect 5244 3516 5252 3524
rect 5404 3516 5412 3524
rect 5596 3516 5604 3524
rect 3548 3496 3556 3504
rect 3628 3496 3636 3504
rect 3644 3496 3652 3504
rect 3676 3496 3684 3504
rect 3740 3496 3748 3504
rect 4204 3496 4212 3504
rect 4300 3496 4308 3504
rect 4396 3496 4404 3504
rect 4460 3496 4468 3504
rect 4908 3496 4916 3504
rect 4988 3496 4996 3504
rect 5116 3496 5124 3504
rect 1740 3476 1748 3484
rect 1772 3476 1780 3484
rect 1980 3476 1988 3484
rect 124 3456 132 3464
rect 380 3456 388 3464
rect 396 3456 404 3464
rect 524 3456 532 3464
rect 620 3456 628 3464
rect 700 3456 708 3464
rect 892 3456 900 3464
rect 1052 3456 1060 3464
rect 1068 3456 1076 3464
rect 1148 3456 1156 3464
rect 1340 3456 1348 3464
rect 1532 3456 1540 3464
rect 1660 3456 1668 3464
rect 1772 3456 1780 3464
rect 1852 3456 1860 3464
rect 1964 3456 1972 3464
rect 2028 3476 2036 3484
rect 2092 3476 2100 3484
rect 2140 3476 2148 3484
rect 2236 3476 2244 3484
rect 2300 3476 2308 3484
rect 2476 3476 2484 3484
rect 2524 3476 2532 3484
rect 2620 3476 2628 3484
rect 2636 3476 2644 3484
rect 2732 3476 2740 3484
rect 2780 3476 2788 3484
rect 2828 3476 2836 3484
rect 2924 3476 2932 3484
rect 2972 3476 2980 3484
rect 3340 3476 3348 3484
rect 3452 3476 3460 3484
rect 3564 3476 3572 3484
rect 3660 3476 3668 3484
rect 3852 3476 3860 3484
rect 3900 3476 3908 3484
rect 3996 3476 4004 3484
rect 4108 3476 4116 3484
rect 4124 3476 4132 3484
rect 4156 3476 4164 3484
rect 4220 3476 4228 3484
rect 4236 3476 4244 3484
rect 4284 3476 4292 3484
rect 4540 3476 4548 3484
rect 4572 3476 4580 3484
rect 4700 3476 4708 3484
rect 4764 3476 4772 3484
rect 4812 3476 4820 3484
rect 4844 3476 4852 3484
rect 4924 3476 4932 3484
rect 5052 3476 5060 3484
rect 5164 3496 5172 3504
rect 5276 3496 5284 3504
rect 5324 3496 5332 3504
rect 5372 3496 5380 3504
rect 5436 3496 5444 3504
rect 5500 3496 5508 3504
rect 5532 3496 5540 3504
rect 5660 3516 5668 3524
rect 5692 3516 5700 3524
rect 5852 3516 5860 3524
rect 5900 3516 5908 3524
rect 6220 3516 6228 3524
rect 5836 3496 5844 3504
rect 5900 3496 5908 3504
rect 5932 3496 5940 3504
rect 6060 3496 6068 3504
rect 5148 3476 5156 3484
rect 5244 3476 5252 3484
rect 5292 3476 5300 3484
rect 5388 3476 5396 3484
rect 5452 3476 5460 3484
rect 5692 3476 5700 3484
rect 5948 3476 5956 3484
rect 6060 3476 6068 3484
rect 6140 3496 6148 3504
rect 6188 3476 6196 3484
rect 6220 3476 6228 3484
rect 2268 3456 2276 3464
rect 2332 3456 2340 3464
rect 2412 3456 2420 3464
rect 2460 3456 2468 3464
rect 2700 3456 2708 3464
rect 2940 3456 2948 3464
rect 3516 3456 3524 3464
rect 3676 3456 3684 3464
rect 3772 3456 3780 3464
rect 3868 3456 3876 3464
rect 4348 3456 4356 3464
rect 4556 3456 4564 3464
rect 4684 3456 4692 3464
rect 4844 3456 4852 3464
rect 4876 3456 4884 3464
rect 5068 3456 5076 3464
rect 5324 3456 5332 3464
rect 5468 3456 5476 3464
rect 5532 3456 5540 3464
rect 5724 3456 5732 3464
rect 5756 3456 5764 3464
rect 5788 3456 5796 3464
rect 5948 3456 5956 3464
rect 412 3436 420 3444
rect 1004 3436 1012 3444
rect 1212 3436 1220 3444
rect 1468 3436 1476 3444
rect 1868 3436 1876 3444
rect 2252 3436 2260 3444
rect 2316 3436 2324 3444
rect 2588 3436 2596 3444
rect 2716 3436 2724 3444
rect 2860 3436 2868 3444
rect 2956 3436 2964 3444
rect 3020 3436 3028 3444
rect 3132 3436 3140 3444
rect 3596 3436 3604 3444
rect 5644 3436 5652 3444
rect 6108 3436 6116 3444
rect 3118 3406 3126 3414
rect 3132 3406 3140 3414
rect 3146 3406 3154 3414
rect 108 3376 116 3384
rect 172 3376 180 3384
rect 188 3376 196 3384
rect 236 3376 244 3384
rect 300 3376 308 3384
rect 348 3376 356 3384
rect 364 3376 372 3384
rect 428 3376 436 3384
rect 700 3376 708 3384
rect 748 3376 756 3384
rect 812 3376 820 3384
rect 860 3376 868 3384
rect 1148 3376 1156 3384
rect 1276 3376 1284 3384
rect 1324 3376 1332 3384
rect 1516 3376 1524 3384
rect 2188 3376 2196 3384
rect 2316 3376 2324 3384
rect 2364 3376 2372 3384
rect 2892 3376 2900 3384
rect 2972 3376 2980 3384
rect 3036 3376 3044 3384
rect 3212 3376 3220 3384
rect 3276 3376 3284 3384
rect 3308 3376 3316 3384
rect 3516 3376 3524 3384
rect 3628 3376 3636 3384
rect 3676 3376 3684 3384
rect 3724 3376 3732 3384
rect 3756 3376 3764 3384
rect 3868 3376 3876 3384
rect 4044 3376 4052 3384
rect 4316 3376 4324 3384
rect 4460 3376 4468 3384
rect 4508 3376 4516 3384
rect 4620 3376 4628 3384
rect 4796 3376 4804 3384
rect 4860 3376 4868 3384
rect 4988 3376 4996 3384
rect 5036 3376 5044 3384
rect 5212 3376 5220 3384
rect 5324 3376 5332 3384
rect 5388 3376 5396 3384
rect 5404 3376 5412 3384
rect 5628 3376 5636 3384
rect 5692 3376 5700 3384
rect 5708 3376 5716 3384
rect 6060 3376 6068 3384
rect 412 3356 420 3364
rect 444 3356 452 3364
rect 588 3356 596 3364
rect 716 3356 724 3364
rect 12 3336 20 3344
rect 156 3336 164 3344
rect 204 3336 212 3344
rect 220 3336 228 3344
rect 252 3336 260 3344
rect 268 3336 276 3344
rect 316 3336 324 3344
rect 396 3336 404 3344
rect 476 3336 484 3344
rect 540 3336 548 3344
rect 604 3336 612 3344
rect 684 3336 692 3344
rect 1052 3356 1060 3364
rect 1116 3356 1124 3364
rect 780 3336 788 3344
rect 828 3336 836 3344
rect 876 3336 884 3344
rect 1036 3336 1044 3344
rect 1228 3356 1236 3364
rect 1372 3356 1380 3364
rect 1612 3356 1620 3364
rect 1868 3356 1876 3364
rect 1980 3356 1988 3364
rect 2556 3356 2564 3364
rect 2572 3356 2580 3364
rect 2844 3356 2852 3364
rect 3052 3356 3060 3364
rect 3196 3356 3204 3364
rect 3324 3356 3332 3364
rect 3740 3356 3748 3364
rect 3852 3356 3860 3364
rect 3932 3356 3940 3364
rect 4060 3356 4068 3364
rect 1244 3336 1252 3344
rect 1292 3336 1300 3344
rect 1340 3336 1348 3344
rect 1388 3336 1396 3344
rect 1436 3336 1444 3344
rect 1452 3336 1460 3344
rect 1548 3336 1556 3344
rect 1644 3336 1652 3344
rect 1660 3336 1668 3344
rect 1724 3336 1732 3344
rect 1788 3336 1796 3344
rect 1868 3336 1876 3344
rect 1932 3336 1940 3344
rect 2156 3336 2164 3344
rect 2252 3336 2260 3344
rect 2540 3336 2548 3344
rect 2764 3336 2772 3344
rect 2796 3336 2804 3344
rect 2828 3336 2836 3344
rect 2908 3336 2916 3344
rect 3004 3336 3012 3344
rect 3228 3336 3236 3344
rect 3292 3336 3300 3344
rect 3340 3336 3348 3344
rect 3372 3336 3380 3344
rect 3468 3336 3476 3344
rect 492 3316 500 3324
rect 556 3316 564 3324
rect 604 3316 612 3324
rect 732 3316 740 3324
rect 940 3316 948 3324
rect 956 3316 964 3324
rect 44 3296 52 3304
rect 172 3296 180 3304
rect 220 3296 228 3304
rect 300 3296 308 3304
rect 348 3296 356 3304
rect 364 3296 372 3304
rect 588 3296 596 3304
rect 652 3296 660 3304
rect 812 3296 820 3304
rect 860 3296 868 3304
rect 908 3296 916 3304
rect 1084 3316 1092 3324
rect 1180 3316 1188 3324
rect 1196 3316 1204 3324
rect 1404 3316 1412 3324
rect 1644 3316 1652 3324
rect 1676 3316 1684 3324
rect 1740 3316 1748 3324
rect 1804 3316 1812 3324
rect 1916 3316 1924 3324
rect 2012 3316 2020 3324
rect 2044 3316 2052 3324
rect 2124 3316 2132 3324
rect 2220 3316 2228 3324
rect 2284 3316 2292 3324
rect 2364 3316 2372 3324
rect 2428 3316 2436 3324
rect 2492 3316 2500 3324
rect 2524 3316 2532 3324
rect 2620 3316 2628 3324
rect 2684 3316 2692 3324
rect 2748 3316 2756 3324
rect 2812 3316 2820 3324
rect 2924 3316 2932 3324
rect 2972 3316 2980 3324
rect 3148 3316 3156 3324
rect 3260 3316 3268 3324
rect 3388 3316 3396 3324
rect 3436 3316 3444 3324
rect 3484 3316 3492 3324
rect 3564 3316 3572 3324
rect 3628 3336 3636 3344
rect 3692 3336 3700 3344
rect 3804 3336 3812 3344
rect 3836 3336 3844 3344
rect 3884 3336 3892 3344
rect 4028 3336 4036 3344
rect 4108 3336 4116 3344
rect 3772 3316 3780 3324
rect 3820 3316 3828 3324
rect 3980 3316 3988 3324
rect 4012 3316 4020 3324
rect 4108 3316 4116 3324
rect 4220 3336 4228 3344
rect 4268 3336 4276 3344
rect 4380 3336 4388 3344
rect 4396 3336 4404 3344
rect 4716 3356 4724 3364
rect 4876 3356 4884 3364
rect 4924 3356 4932 3364
rect 5068 3356 5076 3364
rect 5100 3356 5108 3364
rect 5148 3356 5156 3364
rect 5260 3356 5268 3364
rect 5340 3356 5348 3364
rect 5548 3356 5556 3364
rect 4540 3336 4548 3344
rect 4604 3336 4612 3344
rect 4732 3336 4740 3344
rect 4828 3336 4836 3344
rect 4940 3336 4948 3344
rect 4972 3336 4980 3344
rect 5004 3336 5012 3344
rect 5052 3336 5060 3344
rect 5356 3336 5364 3344
rect 5452 3336 5460 3344
rect 5516 3336 5524 3344
rect 5532 3336 5540 3344
rect 5580 3336 5588 3344
rect 5644 3336 5652 3344
rect 5740 3332 5748 3340
rect 5756 3336 5764 3344
rect 5772 3336 5780 3344
rect 5820 3336 5828 3344
rect 988 3296 996 3304
rect 1276 3296 1284 3304
rect 1324 3296 1332 3304
rect 1372 3296 1380 3304
rect 1436 3296 1444 3304
rect 1772 3296 1780 3304
rect 1884 3296 1892 3304
rect 1932 3296 1940 3304
rect 1964 3296 1972 3304
rect 2044 3296 2052 3304
rect 2156 3296 2164 3304
rect 2188 3296 2196 3304
rect 2204 3296 2212 3304
rect 2316 3296 2324 3304
rect 2380 3296 2388 3304
rect 2444 3296 2452 3304
rect 2508 3296 2516 3304
rect 2636 3296 2644 3304
rect 2700 3296 2708 3304
rect 2716 3296 2724 3304
rect 2780 3296 2788 3304
rect 2988 3296 2996 3304
rect 3036 3296 3044 3304
rect 3164 3296 3172 3304
rect 3260 3296 3268 3304
rect 3452 3296 3460 3304
rect 3580 3296 3588 3304
rect 3644 3296 3652 3304
rect 3676 3296 3684 3304
rect 3724 3296 3732 3304
rect 3788 3296 3796 3304
rect 3996 3296 4004 3304
rect 4076 3296 4084 3304
rect 4236 3296 4244 3304
rect 4428 3296 4436 3304
rect 4492 3316 4500 3324
rect 4556 3316 4564 3324
rect 4844 3316 4852 3324
rect 4892 3316 4900 3324
rect 5100 3316 5108 3324
rect 5116 3316 5124 3324
rect 5180 3316 5188 3324
rect 5228 3316 5236 3324
rect 5292 3316 5300 3324
rect 5436 3316 5444 3324
rect 5452 3316 5460 3324
rect 5500 3316 5508 3324
rect 5596 3316 5604 3324
rect 5660 3316 5668 3324
rect 5788 3316 5796 3324
rect 6140 3356 6148 3364
rect 6220 3356 6228 3364
rect 5852 3336 5860 3344
rect 5964 3336 5972 3344
rect 6012 3336 6020 3344
rect 5900 3316 5908 3324
rect 5980 3316 5988 3324
rect 6124 3336 6132 3344
rect 6188 3316 6196 3324
rect 4588 3296 4596 3304
rect 5020 3296 5028 3304
rect 5052 3296 5060 3304
rect 5212 3296 5220 3304
rect 5324 3296 5332 3304
rect 5468 3296 5476 3304
rect 5580 3296 5588 3304
rect 5820 3296 5828 3304
rect 5916 3296 5924 3304
rect 5932 3296 5940 3304
rect 5980 3296 5988 3304
rect 524 3276 532 3284
rect 1020 3276 1028 3284
rect 1052 3276 1060 3284
rect 1804 3276 1812 3284
rect 2060 3276 2068 3284
rect 2108 3276 2116 3284
rect 2348 3276 2356 3284
rect 2412 3276 2420 3284
rect 2476 3276 2484 3284
rect 2604 3276 2612 3284
rect 2668 3276 2676 3284
rect 2956 3276 2964 3284
rect 3420 3276 3428 3284
rect 3548 3276 3556 3284
rect 3964 3276 3972 3284
rect 4972 3276 4980 3284
rect 5884 3276 5892 3284
rect 460 3256 468 3264
rect 2124 3256 2132 3264
rect 2428 3256 2436 3264
rect 2492 3256 2500 3264
rect 3132 3256 3140 3264
rect 5900 3256 5908 3264
rect 1196 3236 1204 3244
rect 1260 3236 1268 3244
rect 1740 3236 1748 3244
rect 1948 3236 1956 3244
rect 1996 3236 2004 3244
rect 2076 3236 2084 3244
rect 2588 3236 2596 3244
rect 2684 3236 2692 3244
rect 2748 3236 2756 3244
rect 3404 3236 3412 3244
rect 3916 3236 3924 3244
rect 3948 3236 3956 3244
rect 4188 3236 4196 3244
rect 5244 3236 5252 3244
rect 6156 3236 6164 3244
rect 1566 3206 1574 3214
rect 1580 3206 1588 3214
rect 1594 3206 1602 3214
rect 4638 3206 4646 3214
rect 4652 3206 4660 3214
rect 4666 3206 4674 3214
rect 60 3176 68 3184
rect 236 3176 244 3184
rect 316 3176 324 3184
rect 396 3176 404 3184
rect 556 3176 564 3184
rect 892 3176 900 3184
rect 972 3176 980 3184
rect 1180 3176 1188 3184
rect 1804 3176 1812 3184
rect 1964 3176 1972 3184
rect 2252 3176 2260 3184
rect 2348 3176 2356 3184
rect 2732 3176 2740 3184
rect 2860 3176 2868 3184
rect 2940 3176 2948 3184
rect 3036 3176 3044 3184
rect 3164 3176 3172 3184
rect 3212 3176 3220 3184
rect 3308 3176 3316 3184
rect 3372 3176 3380 3184
rect 3500 3176 3508 3184
rect 3708 3176 3716 3184
rect 3884 3176 3892 3184
rect 3980 3176 3988 3184
rect 4572 3176 4580 3184
rect 4716 3176 4724 3184
rect 4860 3176 4868 3184
rect 4924 3176 4932 3184
rect 5260 3176 5268 3184
rect 5468 3176 5476 3184
rect 5548 3176 5556 3184
rect 5644 3176 5652 3184
rect 5708 3176 5716 3184
rect 5836 3176 5844 3184
rect 5916 3176 5924 3184
rect 5964 3176 5972 3184
rect 1148 3156 1156 3164
rect 1324 3156 1332 3164
rect 1868 3156 1876 3164
rect 364 3136 372 3144
rect 524 3136 532 3144
rect 828 3136 836 3144
rect 1132 3136 1140 3144
rect 1308 3136 1316 3144
rect 1516 3136 1524 3144
rect 1532 3136 1540 3144
rect 1644 3136 1652 3144
rect 1996 3136 2004 3144
rect 2092 3136 2100 3144
rect 2108 3136 2116 3144
rect 2636 3136 2644 3144
rect 3260 3156 3268 3164
rect 4172 3156 4180 3164
rect 2876 3136 2884 3144
rect 3052 3136 3060 3144
rect 3292 3136 3300 3144
rect 3420 3136 3428 3144
rect 3532 3136 3540 3144
rect 3596 3136 3604 3144
rect 3628 3136 3636 3144
rect 3788 3136 3796 3144
rect 4092 3136 4100 3144
rect 4156 3136 4164 3144
rect 4540 3136 4548 3144
rect 5372 3136 5380 3144
rect 5660 3136 5668 3144
rect 6188 3136 6196 3144
rect 6236 3136 6244 3144
rect 124 3116 132 3124
rect 172 3116 180 3124
rect 204 3116 212 3124
rect 444 3116 452 3124
rect 588 3116 596 3124
rect 668 3114 676 3122
rect 780 3116 788 3124
rect 796 3116 804 3124
rect 860 3116 868 3124
rect 924 3116 932 3124
rect 1084 3116 1092 3124
rect 1100 3116 1108 3124
rect 1212 3116 1220 3124
rect 1276 3116 1284 3124
rect 1340 3116 1348 3124
rect 1564 3116 1572 3124
rect 1660 3116 1668 3124
rect 1836 3116 1844 3124
rect 1852 3116 1860 3124
rect 2044 3116 2052 3124
rect 2076 3116 2084 3124
rect 2140 3116 2148 3124
rect 2172 3116 2180 3124
rect 2220 3116 2228 3124
rect 2284 3116 2292 3124
rect 2428 3116 2436 3124
rect 2668 3116 2676 3124
rect 2684 3116 2692 3124
rect 2716 3116 2724 3124
rect 2764 3116 2772 3124
rect 2844 3116 2852 3124
rect 2908 3116 2916 3124
rect 3004 3116 3012 3124
rect 3020 3116 3028 3124
rect 3132 3116 3140 3124
rect 3244 3116 3252 3124
rect 3276 3116 3284 3124
rect 3436 3116 3444 3124
rect 3564 3116 3572 3124
rect 3580 3116 3588 3124
rect 3676 3116 3684 3124
rect 380 3096 388 3104
rect 412 3096 420 3104
rect 492 3096 500 3104
rect 556 3096 564 3104
rect 700 3096 708 3104
rect 828 3096 836 3104
rect 892 3096 900 3104
rect 12 3076 20 3084
rect 156 3076 164 3084
rect 204 3076 212 3084
rect 252 3076 260 3084
rect 284 3080 292 3088
rect 332 3076 340 3084
rect 172 3056 180 3064
rect 380 3056 388 3064
rect 412 3056 420 3064
rect 476 3076 484 3084
rect 540 3076 548 3084
rect 652 3076 660 3084
rect 716 3076 724 3084
rect 764 3076 772 3084
rect 812 3076 820 3084
rect 876 3076 884 3084
rect 972 3076 980 3084
rect 1004 3076 1012 3084
rect 1036 3096 1044 3104
rect 1116 3096 1124 3104
rect 1180 3096 1188 3104
rect 1244 3096 1252 3104
rect 1324 3096 1332 3104
rect 1356 3096 1364 3104
rect 1452 3096 1460 3104
rect 1548 3096 1556 3104
rect 1708 3096 1716 3104
rect 1772 3096 1780 3104
rect 1804 3096 1812 3104
rect 1868 3096 1876 3104
rect 1916 3096 1924 3104
rect 2012 3096 2020 3104
rect 2092 3096 2100 3104
rect 2300 3096 2308 3104
rect 2604 3096 2612 3104
rect 2652 3096 2660 3104
rect 2700 3096 2708 3104
rect 2828 3096 2836 3104
rect 2860 3096 2868 3104
rect 2940 3096 2948 3104
rect 1052 3076 1060 3084
rect 1164 3076 1172 3084
rect 1228 3076 1236 3084
rect 1372 3076 1380 3084
rect 1452 3076 1460 3084
rect 1468 3076 1476 3084
rect 1628 3076 1636 3084
rect 1756 3076 1764 3084
rect 1788 3076 1796 3084
rect 1932 3076 1940 3084
rect 2012 3076 2020 3084
rect 2140 3076 2148 3084
rect 2188 3076 2196 3084
rect 2236 3076 2244 3084
rect 2316 3076 2324 3084
rect 2396 3076 2404 3084
rect 2444 3076 2452 3084
rect 2460 3076 2468 3084
rect 2540 3076 2548 3084
rect 620 3056 628 3064
rect 716 3056 724 3064
rect 940 3056 948 3064
rect 972 3056 980 3064
rect 1084 3056 1092 3064
rect 1276 3056 1284 3064
rect 1404 3056 1412 3064
rect 1420 3056 1428 3064
rect 1500 3056 1508 3064
rect 1676 3056 1684 3064
rect 1724 3056 1732 3064
rect 1964 3056 1972 3064
rect 2044 3056 2052 3064
rect 2380 3056 2388 3064
rect 2444 3056 2452 3064
rect 2588 3076 2596 3084
rect 2812 3076 2820 3084
rect 3036 3096 3044 3104
rect 3212 3096 3220 3104
rect 3308 3096 3316 3104
rect 3420 3096 3428 3104
rect 3468 3096 3476 3104
rect 3532 3096 3540 3104
rect 3596 3096 3604 3104
rect 3756 3116 3764 3124
rect 3900 3116 3908 3124
rect 3916 3116 3924 3124
rect 3996 3116 4004 3124
rect 4076 3116 4084 3124
rect 4188 3116 4196 3124
rect 4524 3116 4532 3124
rect 4012 3096 4020 3104
rect 4092 3096 4100 3104
rect 4124 3096 4132 3104
rect 4172 3096 4180 3104
rect 4204 3096 4212 3104
rect 4412 3096 4420 3104
rect 4700 3116 4708 3124
rect 4748 3116 4756 3124
rect 5132 3116 5140 3124
rect 5532 3116 5540 3124
rect 5692 3116 5700 3124
rect 5724 3116 5732 3124
rect 5756 3116 5764 3124
rect 5868 3116 5876 3124
rect 5884 3116 5892 3124
rect 5996 3116 6004 3124
rect 4572 3096 4580 3104
rect 4588 3096 4596 3104
rect 4636 3096 4644 3104
rect 4796 3096 4804 3104
rect 4828 3096 4836 3104
rect 4844 3096 4852 3104
rect 5036 3096 5044 3104
rect 5052 3096 5060 3104
rect 5164 3096 5172 3104
rect 5228 3096 5236 3104
rect 5324 3096 5332 3104
rect 5468 3096 5476 3104
rect 5500 3096 5508 3104
rect 5596 3096 5604 3104
rect 5612 3096 5620 3104
rect 5676 3096 5684 3104
rect 5740 3096 5748 3104
rect 5772 3096 5780 3104
rect 5804 3096 5812 3104
rect 5964 3096 5972 3104
rect 6076 3096 6084 3104
rect 6204 3096 6212 3104
rect 2972 3076 2980 3084
rect 3196 3076 3204 3084
rect 3452 3076 3460 3084
rect 3516 3076 3524 3084
rect 3644 3076 3652 3084
rect 3692 3076 3700 3084
rect 3788 3076 3796 3084
rect 3836 3076 3844 3084
rect 3868 3076 3876 3084
rect 3900 3076 3908 3084
rect 3948 3076 3956 3084
rect 3964 3076 3972 3084
rect 4028 3076 4036 3084
rect 4220 3076 4228 3084
rect 4348 3076 4356 3084
rect 4492 3076 4500 3084
rect 4588 3076 4596 3084
rect 4732 3076 4740 3084
rect 4780 3076 4788 3084
rect 4892 3076 4900 3084
rect 4988 3076 4996 3084
rect 5180 3076 5188 3084
rect 2748 3056 2756 3064
rect 3276 3056 3284 3064
rect 3356 3056 3364 3064
rect 3420 3056 3428 3064
rect 3852 3056 3860 3064
rect 4060 3056 4068 3064
rect 4252 3056 4260 3064
rect 4284 3056 4292 3064
rect 4380 3056 4388 3064
rect 4604 3056 4612 3064
rect 4748 3056 4756 3064
rect 4828 3056 4836 3064
rect 4876 3056 4884 3064
rect 5004 3056 5012 3064
rect 5340 3076 5348 3084
rect 5436 3076 5444 3084
rect 5452 3076 5460 3084
rect 5516 3076 5524 3084
rect 5564 3076 5572 3084
rect 5628 3076 5636 3084
rect 5820 3076 5828 3084
rect 5948 3076 5956 3084
rect 6028 3076 6036 3084
rect 5292 3056 5300 3064
rect 5804 3056 5812 3064
rect 1388 3036 1396 3044
rect 1484 3036 1492 3044
rect 1692 3036 1700 3044
rect 1740 3036 1748 3044
rect 2156 3036 2164 3044
rect 2204 3036 2212 3044
rect 2508 3036 2516 3044
rect 2572 3036 2580 3044
rect 2732 3036 2740 3044
rect 2796 3036 2804 3044
rect 3676 3036 3684 3044
rect 4044 3036 4052 3044
rect 4236 3036 4244 3044
rect 4300 3036 4308 3044
rect 4396 3036 4404 3044
rect 3118 3006 3126 3014
rect 3132 3006 3140 3014
rect 3146 3006 3154 3014
rect 92 2976 100 2984
rect 172 2976 180 2984
rect 268 2976 276 2984
rect 348 2976 356 2984
rect 380 2976 388 2984
rect 412 2976 420 2984
rect 556 2976 564 2984
rect 620 2976 628 2984
rect 716 2976 724 2984
rect 860 2976 868 2984
rect 1004 2976 1012 2984
rect 1148 2976 1156 2984
rect 1340 2976 1348 2984
rect 1612 2976 1620 2984
rect 1676 2976 1684 2984
rect 1836 2976 1844 2984
rect 2268 2976 2276 2984
rect 2556 2976 2564 2984
rect 2812 2976 2820 2984
rect 2876 2976 2884 2984
rect 3036 2976 3044 2984
rect 3100 2976 3108 2984
rect 3244 2976 3252 2984
rect 3324 2976 3332 2984
rect 3420 2976 3428 2984
rect 3516 2976 3524 2984
rect 3708 2976 3716 2984
rect 4092 2976 4100 2984
rect 4156 2976 4164 2984
rect 4572 2976 4580 2984
rect 4716 2976 4724 2984
rect 4732 2976 4740 2984
rect 4892 2976 4900 2984
rect 4940 2976 4948 2984
rect 5068 2976 5076 2984
rect 5436 2976 5444 2984
rect 5516 2976 5524 2984
rect 5644 2976 5652 2984
rect 6012 2976 6020 2984
rect 6092 2976 6100 2984
rect 6124 2976 6132 2984
rect 396 2956 404 2964
rect 524 2956 532 2964
rect 540 2956 548 2964
rect 652 2956 660 2964
rect 780 2956 788 2964
rect 956 2956 964 2964
rect 972 2956 980 2964
rect 988 2956 996 2964
rect 1084 2956 1092 2964
rect 1820 2956 1828 2964
rect 1932 2956 1940 2964
rect 2044 2956 2052 2964
rect 2060 2956 2068 2964
rect 2380 2956 2388 2964
rect 2476 2956 2484 2964
rect 2492 2956 2500 2964
rect 2508 2956 2516 2964
rect 2572 2956 2580 2964
rect 3308 2956 3316 2964
rect 3404 2956 3412 2964
rect 3868 2956 3876 2964
rect 4620 2956 4628 2964
rect 4956 2956 4964 2964
rect 4988 2956 4996 2964
rect 44 2936 52 2944
rect 156 2936 164 2944
rect 204 2936 212 2944
rect 236 2936 244 2944
rect 268 2936 276 2944
rect 300 2936 308 2944
rect 444 2936 452 2944
rect 460 2936 468 2944
rect 588 2936 596 2944
rect 636 2936 644 2944
rect 684 2936 692 2944
rect 732 2936 740 2944
rect 796 2936 804 2944
rect 828 2936 836 2944
rect 860 2936 868 2944
rect 1020 2936 1028 2944
rect 1116 2936 1124 2944
rect 1164 2936 1172 2944
rect 220 2916 228 2924
rect 284 2916 292 2924
rect 316 2916 324 2924
rect 364 2916 372 2924
rect 476 2916 484 2924
rect 748 2916 756 2924
rect 780 2916 788 2924
rect 812 2916 820 2924
rect 908 2916 916 2924
rect 1036 2916 1044 2924
rect 1068 2916 1076 2924
rect 1228 2916 1236 2924
rect 1372 2936 1380 2944
rect 1436 2936 1444 2944
rect 1500 2936 1508 2944
rect 1516 2936 1524 2944
rect 1580 2936 1588 2944
rect 1788 2936 1796 2944
rect 1852 2936 1860 2944
rect 1900 2936 1908 2944
rect 2028 2936 2036 2944
rect 2188 2936 2196 2944
rect 2316 2936 2324 2944
rect 2348 2936 2356 2944
rect 2540 2936 2548 2944
rect 2652 2936 2660 2944
rect 2860 2936 2868 2944
rect 2892 2936 2900 2944
rect 2908 2936 2916 2944
rect 2956 2936 2964 2944
rect 3084 2936 3092 2944
rect 3180 2936 3188 2944
rect 3196 2936 3204 2944
rect 3292 2936 3300 2944
rect 3356 2936 3364 2944
rect 3436 2936 3444 2944
rect 3484 2936 3492 2944
rect 3564 2936 3572 2944
rect 3580 2936 3588 2944
rect 3644 2936 3652 2944
rect 3692 2936 3700 2944
rect 3740 2936 3748 2944
rect 3852 2936 3860 2944
rect 3948 2936 3956 2944
rect 4028 2936 4036 2944
rect 4044 2936 4052 2944
rect 4108 2936 4116 2944
rect 4124 2932 4132 2940
rect 4188 2936 4196 2944
rect 4348 2936 4356 2944
rect 4412 2936 4420 2944
rect 4428 2936 4436 2944
rect 4556 2936 4564 2944
rect 4684 2936 4692 2944
rect 4764 2936 4772 2944
rect 4812 2936 4820 2944
rect 1420 2916 1428 2924
rect 1468 2916 1476 2924
rect 1484 2916 1492 2924
rect 1532 2916 1540 2924
rect 1644 2916 1652 2924
rect 1724 2916 1732 2924
rect 1788 2916 1796 2924
rect 1868 2916 1876 2924
rect 1884 2916 1892 2924
rect 1980 2916 1988 2924
rect 2012 2916 2020 2924
rect 2108 2916 2116 2924
rect 2172 2916 2180 2924
rect 2268 2916 2276 2924
rect 2300 2916 2308 2924
rect 2332 2916 2340 2924
rect 2412 2916 2420 2924
rect 2524 2916 2532 2924
rect 2620 2916 2628 2924
rect 2732 2916 2740 2924
rect 2764 2916 2772 2924
rect 2812 2916 2820 2924
rect 2908 2916 2916 2924
rect 3004 2916 3012 2924
rect 3068 2916 3076 2924
rect 3212 2916 3220 2924
rect 3340 2916 3348 2924
rect 3404 2916 3412 2924
rect 3484 2916 3492 2924
rect 3596 2916 3604 2924
rect 3820 2916 3828 2924
rect 3836 2916 3844 2924
rect 4012 2916 4020 2924
rect 4060 2916 4068 2924
rect 4204 2916 4212 2924
rect 4252 2916 4260 2924
rect 4300 2916 4308 2924
rect 4380 2916 4388 2924
rect 4460 2916 4468 2924
rect 4492 2916 4500 2924
rect 4540 2916 4548 2924
rect 4924 2936 4932 2944
rect 5100 2936 5108 2944
rect 5132 2936 5140 2944
rect 5164 2936 5172 2944
rect 5212 2956 5220 2964
rect 5468 2956 5476 2964
rect 5740 2956 5748 2964
rect 5868 2956 5876 2964
rect 5900 2956 5908 2964
rect 5932 2956 5940 2964
rect 5372 2936 5380 2944
rect 5452 2936 5460 2944
rect 5532 2936 5540 2944
rect 5596 2936 5604 2944
rect 5612 2936 5620 2944
rect 5740 2936 5748 2944
rect 5772 2936 5780 2944
rect 5852 2936 5860 2944
rect 6060 2936 6068 2944
rect 6108 2936 6116 2944
rect 6156 2936 6164 2944
rect 5036 2916 5044 2924
rect 5148 2916 5156 2924
rect 5244 2916 5252 2924
rect 5356 2916 5364 2924
rect 5548 2916 5556 2924
rect 5676 2916 5684 2924
rect 5724 2916 5732 2924
rect 5788 2916 5796 2924
rect 5804 2916 5812 2924
rect 5836 2916 5844 2924
rect 5900 2916 5908 2924
rect 5964 2916 5972 2924
rect 6060 2916 6068 2924
rect 6188 2916 6196 2924
rect 12 2896 20 2904
rect 172 2896 180 2904
rect 540 2896 548 2904
rect 604 2896 612 2904
rect 716 2896 724 2904
rect 892 2896 900 2904
rect 1068 2896 1076 2904
rect 1148 2896 1156 2904
rect 1228 2896 1236 2904
rect 1388 2896 1396 2904
rect 1452 2896 1460 2904
rect 1612 2896 1620 2904
rect 1676 2896 1684 2904
rect 1740 2896 1748 2904
rect 1804 2896 1812 2904
rect 1948 2896 1956 2904
rect 2124 2896 2132 2904
rect 2140 2896 2148 2904
rect 2252 2896 2260 2904
rect 2268 2896 2276 2904
rect 2396 2896 2404 2904
rect 2588 2896 2596 2904
rect 2700 2896 2708 2904
rect 2716 2896 2724 2904
rect 2828 2896 2836 2904
rect 2924 2896 2932 2904
rect 3004 2896 3012 2904
rect 3148 2896 3156 2904
rect 3260 2896 3268 2904
rect 3292 2896 3300 2904
rect 3388 2896 3396 2904
rect 3484 2896 3492 2904
rect 3516 2896 3524 2904
rect 3532 2896 3540 2904
rect 3724 2896 3732 2904
rect 3980 2896 3988 2904
rect 4092 2896 4100 2904
rect 4220 2896 4228 2904
rect 4300 2896 4308 2904
rect 4412 2896 4420 2904
rect 4460 2896 4468 2904
rect 4476 2896 4484 2904
rect 4716 2896 4724 2904
rect 4780 2896 4788 2904
rect 5052 2896 5060 2904
rect 5068 2896 5076 2904
rect 5100 2896 5108 2904
rect 5404 2896 5412 2904
rect 5420 2896 5428 2904
rect 5564 2896 5572 2904
rect 5644 2896 5652 2904
rect 5660 2896 5668 2904
rect 5996 2896 6004 2904
rect 6012 2896 6020 2904
rect 6076 2896 6084 2904
rect 6124 2896 6132 2904
rect 6172 2896 6180 2904
rect 412 2876 420 2884
rect 924 2876 932 2884
rect 1708 2876 1716 2884
rect 1772 2876 1780 2884
rect 1932 2876 1940 2884
rect 1964 2876 1972 2884
rect 2092 2876 2100 2884
rect 2428 2876 2436 2884
rect 2460 2876 2468 2884
rect 2668 2876 2676 2884
rect 2796 2876 2804 2884
rect 2988 2876 2996 2884
rect 3564 2876 3572 2884
rect 4252 2876 4260 2884
rect 4268 2876 4276 2884
rect 4508 2876 4516 2884
rect 5020 2876 5028 2884
rect 5692 2876 5700 2884
rect 6188 2876 6196 2884
rect 668 2856 676 2864
rect 1100 2856 1108 2864
rect 5676 2856 5684 2864
rect 508 2836 516 2844
rect 908 2836 916 2844
rect 1004 2836 1012 2844
rect 1036 2836 1044 2844
rect 1132 2836 1140 2844
rect 1420 2836 1428 2844
rect 1724 2836 1732 2844
rect 1996 2836 2004 2844
rect 2076 2836 2084 2844
rect 2172 2836 2180 2844
rect 2380 2836 2388 2844
rect 2412 2836 2420 2844
rect 2620 2836 2628 2844
rect 3004 2836 3012 2844
rect 3596 2836 3604 2844
rect 3948 2836 3956 2844
rect 4252 2836 4260 2844
rect 4380 2836 4388 2844
rect 4492 2836 4500 2844
rect 4940 2836 4948 2844
rect 4972 2836 4980 2844
rect 5004 2836 5012 2844
rect 5292 2836 5300 2844
rect 5580 2836 5588 2844
rect 5900 2836 5908 2844
rect 5964 2836 5972 2844
rect 6220 2836 6228 2844
rect 1566 2806 1574 2814
rect 1580 2806 1588 2814
rect 1594 2806 1602 2814
rect 4638 2806 4646 2814
rect 4652 2806 4660 2814
rect 4666 2806 4674 2814
rect 44 2776 52 2784
rect 92 2776 100 2784
rect 188 2776 196 2784
rect 236 2776 244 2784
rect 636 2776 644 2784
rect 1276 2776 1284 2784
rect 1836 2776 1844 2784
rect 2108 2776 2116 2784
rect 2140 2776 2148 2784
rect 2748 2776 2756 2784
rect 2844 2776 2852 2784
rect 2924 2776 2932 2784
rect 2988 2776 2996 2784
rect 3100 2776 3108 2784
rect 3196 2776 3204 2784
rect 3548 2776 3556 2784
rect 3884 2776 3892 2784
rect 3996 2776 4004 2784
rect 4236 2776 4244 2784
rect 4476 2776 4484 2784
rect 4588 2776 4596 2784
rect 5148 2776 5156 2784
rect 5212 2776 5220 2784
rect 5356 2776 5364 2784
rect 5484 2776 5492 2784
rect 5756 2776 5764 2784
rect 5932 2776 5940 2784
rect 6220 2776 6228 2784
rect 476 2756 484 2764
rect 764 2756 772 2764
rect 2428 2756 2436 2764
rect 3820 2756 3828 2764
rect 5516 2756 5524 2764
rect 748 2736 756 2744
rect 892 2736 900 2744
rect 2092 2736 2100 2744
rect 2236 2736 2244 2744
rect 2284 2736 2292 2744
rect 2412 2736 2420 2744
rect 2908 2736 2916 2744
rect 2972 2736 2980 2744
rect 3084 2736 3092 2744
rect 3196 2736 3204 2744
rect 3804 2736 3812 2744
rect 3868 2736 3876 2744
rect 3964 2736 3972 2744
rect 3980 2736 3988 2744
rect 4044 2736 4052 2744
rect 4220 2736 4228 2744
rect 4428 2736 4436 2744
rect 4492 2736 4500 2744
rect 4508 2736 4516 2744
rect 108 2716 116 2724
rect 284 2716 292 2724
rect 444 2716 452 2724
rect 540 2716 548 2724
rect 604 2716 612 2724
rect 652 2716 660 2724
rect 716 2716 724 2724
rect 780 2716 788 2724
rect 860 2716 868 2724
rect 1004 2716 1012 2724
rect 1084 2716 1092 2724
rect 1100 2716 1108 2724
rect 1404 2716 1412 2724
rect 1468 2716 1476 2724
rect 1516 2716 1524 2724
rect 1532 2716 1540 2724
rect 1644 2716 1652 2724
rect 1676 2716 1684 2724
rect 1740 2716 1748 2724
rect 2124 2716 2132 2724
rect 2204 2716 2212 2724
rect 2316 2716 2324 2724
rect 2444 2716 2452 2724
rect 2588 2716 2596 2724
rect 2716 2716 2724 2724
rect 2796 2716 2804 2724
rect 2812 2716 2820 2724
rect 2876 2716 2884 2724
rect 2940 2716 2948 2724
rect 2988 2716 2996 2724
rect 3020 2716 3028 2724
rect 3052 2716 3060 2724
rect 3100 2716 3108 2724
rect 3180 2716 3188 2724
rect 3244 2716 3252 2724
rect 3292 2716 3300 2724
rect 3388 2716 3396 2724
rect 12 2696 20 2704
rect 60 2696 68 2704
rect 156 2696 164 2704
rect 204 2696 212 2704
rect 316 2696 324 2704
rect 364 2696 372 2704
rect 396 2696 404 2704
rect 572 2696 580 2704
rect 652 2696 660 2704
rect 684 2696 692 2704
rect 764 2696 772 2704
rect 796 2696 804 2704
rect 908 2696 916 2704
rect 940 2696 948 2704
rect 44 2676 52 2684
rect 140 2676 148 2684
rect 252 2676 260 2684
rect 284 2676 292 2684
rect 412 2676 420 2684
rect 492 2676 500 2684
rect 508 2680 516 2688
rect 556 2676 564 2684
rect 620 2676 628 2684
rect 668 2676 676 2684
rect 812 2676 820 2684
rect 892 2676 900 2684
rect 956 2676 964 2684
rect 1052 2696 1060 2704
rect 1132 2696 1140 2704
rect 1164 2696 1172 2704
rect 1228 2696 1236 2704
rect 1260 2696 1268 2704
rect 1292 2696 1300 2704
rect 1324 2696 1332 2704
rect 1436 2696 1444 2704
rect 1564 2696 1572 2704
rect 1692 2696 1700 2704
rect 1788 2696 1796 2704
rect 1852 2696 1860 2704
rect 1980 2696 1988 2704
rect 2028 2696 2036 2704
rect 2108 2696 2116 2704
rect 2188 2696 2196 2704
rect 2220 2696 2228 2704
rect 2300 2696 2308 2704
rect 2332 2696 2340 2704
rect 2428 2696 2436 2704
rect 2460 2696 2468 2704
rect 2572 2696 2580 2704
rect 2604 2696 2612 2704
rect 2668 2696 2676 2704
rect 2700 2696 2708 2704
rect 2748 2696 2756 2704
rect 1052 2676 1060 2684
rect 1148 2676 1156 2684
rect 1180 2676 1188 2684
rect 1212 2676 1220 2684
rect 1228 2676 1236 2684
rect 1308 2676 1316 2684
rect 1372 2676 1380 2684
rect 1420 2676 1428 2684
rect 1484 2676 1492 2684
rect 1548 2676 1556 2684
rect 1580 2676 1588 2684
rect 1676 2676 1684 2684
rect 1692 2676 1700 2684
rect 1884 2676 1892 2684
rect 1964 2676 1972 2684
rect 2060 2676 2068 2684
rect 2172 2676 2180 2684
rect 2252 2676 2260 2684
rect 2284 2676 2292 2684
rect 2348 2676 2356 2684
rect 2476 2676 2484 2684
rect 2524 2676 2532 2684
rect 2684 2676 2692 2684
rect 2780 2696 2788 2704
rect 2844 2696 2852 2704
rect 2924 2696 2932 2704
rect 2988 2696 2996 2704
rect 3100 2696 3108 2704
rect 3196 2696 3204 2704
rect 3356 2696 3364 2704
rect 3436 2716 3444 2724
rect 3516 2716 3524 2724
rect 3772 2716 3780 2724
rect 3836 2716 3844 2724
rect 3948 2716 3956 2724
rect 4012 2716 4020 2724
rect 4060 2716 4068 2724
rect 4108 2716 4116 2724
rect 4172 2716 4180 2724
rect 4252 2716 4260 2724
rect 4396 2716 4404 2724
rect 4460 2716 4468 2724
rect 4524 2716 4532 2724
rect 4572 2736 4580 2744
rect 5132 2736 5140 2744
rect 5196 2736 5204 2744
rect 5244 2736 5252 2744
rect 5308 2736 5316 2744
rect 5500 2736 5508 2744
rect 5740 2736 5748 2744
rect 4796 2716 4804 2724
rect 4860 2716 4868 2724
rect 3468 2696 3476 2704
rect 3644 2696 3652 2704
rect 3740 2696 3748 2704
rect 3772 2696 3780 2704
rect 3820 2696 3828 2704
rect 3884 2696 3892 2704
rect 3964 2696 3972 2704
rect 4028 2696 4036 2704
rect 4092 2696 4100 2704
rect 4124 2696 4132 2704
rect 4188 2696 4196 2704
rect 4236 2696 4244 2704
rect 4300 2696 4308 2704
rect 4332 2696 4340 2704
rect 4364 2696 4372 2704
rect 4428 2696 4436 2704
rect 4508 2696 4516 2704
rect 4556 2696 4564 2704
rect 4604 2696 4612 2704
rect 4700 2696 4708 2704
rect 4828 2696 4836 2704
rect 4956 2716 4964 2724
rect 5036 2716 5044 2724
rect 5068 2716 5076 2724
rect 5084 2716 5092 2724
rect 5164 2716 5172 2724
rect 5372 2716 5380 2724
rect 5468 2716 5476 2724
rect 5532 2716 5540 2724
rect 5564 2716 5572 2724
rect 5660 2716 5668 2724
rect 5708 2716 5716 2724
rect 5772 2716 5780 2724
rect 5900 2716 5908 2724
rect 6012 2716 6020 2724
rect 6076 2716 6084 2724
rect 6124 2716 6132 2724
rect 5068 2696 5076 2704
rect 5148 2696 5156 2704
rect 5212 2696 5220 2704
rect 5292 2696 5300 2704
rect 5340 2696 5348 2704
rect 5372 2696 5380 2704
rect 5484 2696 5492 2704
rect 5564 2696 5572 2704
rect 5724 2696 5732 2704
rect 5820 2696 5828 2704
rect 5900 2696 5908 2704
rect 6012 2696 6020 2704
rect 6044 2696 6052 2704
rect 6172 2696 6180 2704
rect 2780 2676 2788 2684
rect 2828 2676 2836 2684
rect 3020 2676 3028 2684
rect 3276 2676 3284 2684
rect 3324 2676 3332 2684
rect 3340 2676 3348 2684
rect 3468 2676 3476 2684
rect 3516 2676 3524 2684
rect 3532 2676 3540 2684
rect 3724 2676 3732 2684
rect 4076 2676 4084 2684
rect 4108 2676 4116 2684
rect 4172 2676 4180 2684
rect 4284 2676 4292 2684
rect 4316 2676 4324 2684
rect 4348 2676 4356 2684
rect 4412 2676 4420 2684
rect 364 2656 372 2664
rect 460 2656 468 2664
rect 716 2656 724 2664
rect 908 2656 916 2664
rect 924 2656 932 2664
rect 988 2656 996 2664
rect 1068 2656 1076 2664
rect 1356 2656 1364 2664
rect 1756 2656 1764 2664
rect 1884 2656 1892 2664
rect 1900 2656 1908 2664
rect 2060 2656 2068 2664
rect 2140 2656 2148 2664
rect 2380 2656 2388 2664
rect 2508 2656 2516 2664
rect 2588 2656 2596 2664
rect 2620 2656 2628 2664
rect 3596 2656 3604 2664
rect 3660 2656 3668 2664
rect 3916 2656 3924 2664
rect 4396 2656 4404 2664
rect 4652 2656 4660 2664
rect 4748 2676 4756 2684
rect 4764 2676 4772 2684
rect 4812 2676 4820 2684
rect 4908 2676 4916 2684
rect 4924 2676 4932 2684
rect 4988 2676 4996 2684
rect 5036 2676 5044 2684
rect 5388 2676 5396 2684
rect 5436 2676 5444 2684
rect 5580 2676 5588 2684
rect 5628 2676 5636 2684
rect 5692 2676 5700 2684
rect 5772 2676 5780 2684
rect 5900 2676 5908 2684
rect 5964 2676 5972 2684
rect 6028 2676 6036 2684
rect 6108 2676 6116 2684
rect 6156 2676 6164 2684
rect 6204 2676 6212 2684
rect 4748 2656 4756 2664
rect 4972 2656 4980 2664
rect 5100 2656 5108 2664
rect 5244 2656 5252 2664
rect 5596 2656 5604 2664
rect 5644 2656 5652 2664
rect 5836 2656 5844 2664
rect 5916 2656 5924 2664
rect 5948 2656 5956 2664
rect 6140 2656 6148 2664
rect 6236 2656 6244 2664
rect 124 2636 132 2644
rect 188 2636 196 2644
rect 236 2636 244 2644
rect 268 2636 276 2644
rect 380 2636 388 2644
rect 444 2636 452 2644
rect 604 2636 612 2644
rect 828 2636 836 2644
rect 972 2636 980 2644
rect 1020 2636 1028 2644
rect 1100 2636 1108 2644
rect 1196 2636 1204 2644
rect 1340 2636 1348 2644
rect 1404 2636 1412 2644
rect 1468 2636 1476 2644
rect 1516 2636 1524 2644
rect 1740 2636 1748 2644
rect 1868 2636 1876 2644
rect 1948 2636 1956 2644
rect 2012 2636 2020 2644
rect 2364 2636 2372 2644
rect 3260 2636 3268 2644
rect 3308 2636 3316 2644
rect 4780 2636 4788 2644
rect 4956 2636 4964 2644
rect 5436 2636 5444 2644
rect 5484 2636 5492 2644
rect 5660 2636 5668 2644
rect 5852 2636 5860 2644
rect 6076 2636 6084 2644
rect 3118 2606 3126 2614
rect 3132 2606 3140 2614
rect 3146 2606 3154 2614
rect 92 2576 100 2584
rect 204 2576 212 2584
rect 252 2576 260 2584
rect 652 2576 660 2584
rect 716 2576 724 2584
rect 828 2576 836 2584
rect 1068 2576 1076 2584
rect 1628 2576 1636 2584
rect 1788 2576 1796 2584
rect 2044 2576 2052 2584
rect 2636 2576 2644 2584
rect 2780 2576 2788 2584
rect 3036 2576 3044 2584
rect 3212 2576 3220 2584
rect 3388 2576 3396 2584
rect 3468 2576 3476 2584
rect 3548 2576 3556 2584
rect 3628 2576 3636 2584
rect 3932 2576 3940 2584
rect 4140 2576 4148 2584
rect 4188 2576 4196 2584
rect 4428 2576 4436 2584
rect 4508 2576 4516 2584
rect 4540 2576 4548 2584
rect 4876 2576 4884 2584
rect 5020 2576 5028 2584
rect 5548 2576 5556 2584
rect 5740 2576 5748 2584
rect 5756 2576 5764 2584
rect 5804 2576 5812 2584
rect 6156 2576 6164 2584
rect 332 2556 340 2564
rect 348 2556 356 2564
rect 572 2556 580 2564
rect 636 2556 644 2564
rect 908 2556 916 2564
rect 1100 2556 1108 2564
rect 1148 2556 1156 2564
rect 1516 2556 1524 2564
rect 1772 2556 1780 2564
rect 1804 2556 1812 2564
rect 1948 2556 1956 2564
rect 348 2536 356 2544
rect 508 2536 516 2544
rect 556 2536 564 2544
rect 620 2536 628 2544
rect 668 2536 676 2544
rect 748 2536 756 2544
rect 860 2536 868 2544
rect 972 2536 980 2544
rect 1052 2536 1060 2544
rect 1132 2536 1140 2544
rect 1276 2536 1284 2544
rect 1292 2536 1300 2544
rect 1388 2536 1396 2544
rect 1484 2536 1492 2544
rect 1532 2536 1540 2544
rect 1612 2536 1620 2544
rect 1820 2536 1828 2544
rect 1980 2536 1988 2544
rect 1996 2536 2004 2544
rect 2076 2556 2084 2564
rect 2364 2556 2372 2564
rect 2460 2556 2468 2564
rect 2796 2556 2804 2564
rect 3020 2556 3028 2564
rect 3196 2556 3204 2564
rect 3644 2556 3652 2564
rect 3772 2556 3780 2564
rect 4076 2556 4084 2564
rect 4092 2556 4100 2564
rect 4204 2556 4212 2564
rect 4380 2556 4388 2564
rect 4796 2556 4804 2564
rect 2108 2536 2116 2544
rect 2300 2536 2308 2544
rect 2380 2536 2388 2544
rect 2652 2536 2660 2544
rect 2732 2536 2740 2544
rect 3116 2536 3124 2544
rect 3228 2536 3236 2544
rect 3372 2536 3380 2544
rect 3420 2536 3428 2544
rect 3436 2536 3444 2544
rect 3484 2536 3492 2544
rect 3548 2536 3556 2544
rect 3580 2536 3588 2544
rect 3660 2536 3668 2544
rect 3692 2536 3700 2544
rect 3724 2536 3732 2544
rect 3756 2536 3764 2544
rect 3804 2536 3812 2544
rect 3932 2536 3940 2544
rect 3964 2536 3972 2544
rect 3996 2536 4004 2544
rect 4060 2536 4068 2544
rect 4284 2536 4292 2544
rect 4332 2536 4340 2544
rect 4396 2536 4404 2544
rect 4412 2536 4420 2544
rect 4476 2536 4484 2544
rect 4524 2536 4532 2544
rect 4588 2536 4596 2544
rect 4652 2536 4660 2544
rect 12 2516 20 2524
rect 60 2516 68 2524
rect 124 2516 132 2524
rect 172 2516 180 2524
rect 220 2516 228 2524
rect 300 2516 308 2524
rect 380 2516 388 2524
rect 396 2516 404 2524
rect 460 2516 468 2524
rect 524 2516 532 2524
rect 556 2516 564 2524
rect 604 2516 612 2524
rect 684 2516 692 2524
rect 764 2516 772 2524
rect 828 2516 836 2524
rect 860 2516 868 2524
rect 924 2516 932 2524
rect 956 2516 964 2524
rect 1436 2516 1444 2524
rect 1532 2516 1540 2524
rect 1548 2516 1556 2524
rect 1660 2516 1668 2524
rect 1740 2516 1748 2524
rect 1804 2516 1812 2524
rect 1900 2516 1908 2524
rect 1996 2516 2004 2524
rect 2012 2516 2020 2524
rect 2124 2516 2132 2524
rect 2204 2516 2212 2524
rect 2252 2516 2260 2524
rect 2316 2516 2324 2524
rect 2332 2516 2340 2524
rect 2412 2516 2420 2524
rect 2444 2516 2452 2524
rect 2508 2516 2516 2524
rect 2572 2516 2580 2524
rect 2700 2516 2708 2524
rect 2844 2516 2852 2524
rect 2876 2516 2884 2524
rect 2924 2516 2932 2524
rect 2972 2516 2980 2524
rect 3068 2516 3076 2524
rect 3148 2516 3156 2524
rect 3260 2516 3268 2524
rect 3308 2516 3316 2524
rect 3388 2516 3396 2524
rect 3500 2516 3508 2524
rect 3532 2516 3540 2524
rect 108 2496 116 2504
rect 316 2496 324 2504
rect 412 2496 420 2504
rect 476 2496 484 2504
rect 572 2496 580 2504
rect 780 2496 788 2504
rect 844 2496 852 2504
rect 924 2496 932 2504
rect 1036 2496 1044 2504
rect 1084 2496 1092 2504
rect 1100 2496 1108 2504
rect 1436 2496 1444 2504
rect 1580 2496 1588 2504
rect 1692 2496 1700 2504
rect 1708 2496 1716 2504
rect 1868 2496 1876 2504
rect 1884 2496 1892 2504
rect 2156 2496 2164 2504
rect 2220 2496 2228 2504
rect 2236 2496 2244 2504
rect 2348 2496 2356 2504
rect 2396 2496 2404 2504
rect 2476 2496 2484 2504
rect 2556 2496 2564 2504
rect 2652 2496 2660 2504
rect 2668 2496 2676 2504
rect 2700 2496 2708 2504
rect 2828 2496 2836 2504
rect 2940 2496 2948 2504
rect 3132 2496 3140 2504
rect 3292 2496 3300 2504
rect 3324 2496 3332 2504
rect 3388 2496 3396 2504
rect 3468 2496 3476 2504
rect 3532 2496 3540 2504
rect 3596 2516 3604 2524
rect 3676 2496 3684 2504
rect 3740 2516 3748 2524
rect 3788 2516 3796 2524
rect 3884 2516 3892 2524
rect 3916 2516 3924 2524
rect 3980 2516 3988 2524
rect 4012 2516 4020 2524
rect 4140 2516 4148 2524
rect 4252 2516 4260 2524
rect 4300 2516 4308 2524
rect 4460 2516 4468 2524
rect 3708 2496 3716 2504
rect 3836 2496 3844 2504
rect 3900 2496 3908 2504
rect 4044 2496 4052 2504
rect 4124 2496 4132 2504
rect 4268 2496 4276 2504
rect 4316 2496 4324 2504
rect 4428 2496 4436 2504
rect 4572 2516 4580 2524
rect 4732 2516 4740 2524
rect 4764 2516 4772 2524
rect 5004 2536 5012 2544
rect 5052 2556 5060 2564
rect 5084 2556 5092 2564
rect 5148 2556 5156 2564
rect 5292 2556 5300 2564
rect 5852 2556 5860 2564
rect 5212 2536 5220 2544
rect 5372 2536 5380 2544
rect 5436 2536 5444 2544
rect 5468 2536 5476 2544
rect 5580 2536 5588 2544
rect 5596 2536 5604 2544
rect 5708 2536 5716 2544
rect 5788 2536 5796 2544
rect 5836 2536 5844 2544
rect 5884 2536 5892 2544
rect 5932 2536 5940 2544
rect 6028 2536 6036 2544
rect 6108 2536 6116 2544
rect 4588 2496 4596 2504
rect 4764 2496 4772 2504
rect 4812 2496 4820 2504
rect 140 2476 148 2484
rect 284 2476 292 2484
rect 444 2476 452 2484
rect 748 2476 756 2484
rect 812 2476 820 2484
rect 1228 2476 1236 2484
rect 1356 2476 1364 2484
rect 1420 2476 1428 2484
rect 1916 2476 1924 2484
rect 2188 2476 2196 2484
rect 2204 2476 2212 2484
rect 1004 2456 1012 2464
rect 2124 2456 2132 2464
rect 2268 2476 2276 2484
rect 2428 2476 2436 2484
rect 2524 2476 2532 2484
rect 2572 2476 2580 2484
rect 2908 2476 2916 2484
rect 2988 2476 2996 2484
rect 3116 2476 3124 2484
rect 3164 2476 3172 2484
rect 3868 2476 3876 2484
rect 4236 2476 4244 2484
rect 4636 2476 4644 2484
rect 4796 2476 4804 2484
rect 4940 2516 4948 2524
rect 4988 2516 4996 2524
rect 5132 2516 5140 2524
rect 5244 2516 5252 2524
rect 5324 2516 5332 2524
rect 5388 2516 5396 2524
rect 5516 2516 5524 2524
rect 6028 2516 6036 2524
rect 6076 2516 6084 2524
rect 6188 2516 6196 2524
rect 4876 2496 4884 2504
rect 4924 2496 4932 2504
rect 5164 2496 5172 2504
rect 5196 2496 5204 2504
rect 5276 2496 5284 2504
rect 5420 2496 5428 2504
rect 5468 2496 5476 2504
rect 5532 2496 5540 2504
rect 5548 2496 5556 2504
rect 5740 2496 5748 2504
rect 5788 2496 5796 2504
rect 5916 2496 5924 2504
rect 6044 2496 6052 2504
rect 6156 2496 6164 2504
rect 4844 2476 4852 2484
rect 4860 2476 4868 2484
rect 4956 2476 4964 2484
rect 5244 2476 5252 2484
rect 5340 2476 5348 2484
rect 5500 2476 5508 2484
rect 5660 2476 5668 2484
rect 6204 2476 6212 2484
rect 3820 2456 3828 2464
rect 3884 2456 3892 2464
rect 5516 2456 5524 2464
rect 44 2436 52 2444
rect 92 2436 100 2444
rect 156 2436 164 2444
rect 204 2436 212 2444
rect 252 2436 260 2444
rect 300 2436 308 2444
rect 460 2436 468 2444
rect 956 2436 964 2444
rect 1436 2436 1444 2444
rect 1660 2436 1668 2444
rect 1724 2436 1732 2444
rect 1836 2436 1844 2444
rect 1900 2436 1908 2444
rect 1948 2436 1956 2444
rect 2172 2436 2180 2444
rect 2508 2436 2516 2444
rect 2572 2436 2580 2444
rect 2844 2436 2852 2444
rect 2924 2436 2932 2444
rect 2972 2436 2980 2444
rect 4012 2436 4020 2444
rect 4252 2436 4260 2444
rect 4732 2436 4740 2444
rect 4940 2436 4948 2444
rect 5900 2436 5908 2444
rect 5964 2436 5972 2444
rect 6188 2436 6196 2444
rect 1566 2406 1574 2414
rect 1580 2406 1588 2414
rect 1594 2406 1602 2414
rect 4638 2406 4646 2414
rect 4652 2406 4660 2414
rect 4666 2406 4674 2414
rect 508 2376 516 2384
rect 1068 2376 1076 2384
rect 2476 2376 2484 2384
rect 2588 2376 2596 2384
rect 2668 2376 2676 2384
rect 2764 2376 2772 2384
rect 2940 2376 2948 2384
rect 2972 2376 2980 2384
rect 3836 2376 3844 2384
rect 4124 2376 4132 2384
rect 4812 2376 4820 2384
rect 5388 2376 5396 2384
rect 5660 2376 5668 2384
rect 5820 2376 5828 2384
rect 6076 2376 6084 2384
rect 3340 2356 3348 2364
rect 5548 2356 5556 2364
rect 5868 2356 5876 2364
rect 92 2336 100 2344
rect 268 2336 276 2344
rect 316 2336 324 2344
rect 652 2336 660 2344
rect 972 2336 980 2344
rect 1180 2336 1188 2344
rect 1340 2336 1348 2344
rect 1708 2336 1716 2344
rect 1852 2336 1860 2344
rect 1900 2336 1908 2344
rect 1964 2336 1972 2344
rect 2316 2336 2324 2344
rect 2364 2336 2372 2344
rect 2396 2336 2404 2344
rect 2460 2336 2468 2344
rect 2572 2336 2580 2344
rect 2636 2336 2644 2344
rect 2684 2336 2692 2344
rect 2716 2336 2724 2344
rect 2748 2336 2756 2344
rect 2812 2336 2820 2344
rect 2844 2336 2852 2344
rect 2860 2336 2868 2344
rect 2892 2336 2900 2344
rect 3324 2336 3332 2344
rect 3644 2336 3652 2344
rect 3772 2336 3780 2344
rect 3820 2336 3828 2344
rect 3932 2336 3940 2344
rect 3964 2336 3972 2344
rect 4284 2336 4292 2344
rect 5212 2336 5220 2344
rect 5404 2336 5412 2344
rect 5564 2336 5572 2344
rect 5804 2336 5812 2344
rect 5868 2336 5876 2344
rect 5916 2336 5924 2344
rect 6028 2336 6036 2344
rect 12 2316 20 2324
rect 60 2316 68 2324
rect 188 2316 196 2324
rect 284 2316 292 2324
rect 348 2316 356 2324
rect 684 2316 692 2324
rect 748 2316 756 2324
rect 188 2296 196 2304
rect 220 2296 228 2304
rect 332 2296 340 2304
rect 364 2296 372 2304
rect 428 2296 436 2304
rect 492 2296 500 2304
rect 572 2296 580 2304
rect 652 2296 660 2304
rect 716 2296 724 2304
rect 828 2316 836 2324
rect 860 2316 868 2324
rect 940 2316 948 2324
rect 1004 2316 1012 2324
rect 1100 2316 1108 2324
rect 1212 2316 1220 2324
rect 1372 2316 1380 2324
rect 1452 2316 1460 2324
rect 1516 2316 1524 2324
rect 1676 2316 1684 2324
rect 1740 2316 1748 2324
rect 1820 2316 1828 2324
rect 1932 2316 1940 2324
rect 1948 2316 1956 2324
rect 1996 2316 2004 2324
rect 2012 2316 2020 2324
rect 2060 2316 2068 2324
rect 2236 2316 2244 2324
rect 2364 2316 2372 2324
rect 2428 2316 2436 2324
rect 2604 2316 2612 2324
rect 2716 2316 2724 2324
rect 2892 2316 2900 2324
rect 828 2296 836 2304
rect 908 2296 916 2304
rect 988 2296 996 2304
rect 1020 2296 1028 2304
rect 1084 2296 1092 2304
rect 1132 2296 1140 2304
rect 1196 2296 1204 2304
rect 1292 2296 1300 2304
rect 1356 2296 1364 2304
rect 1452 2296 1460 2304
rect 1484 2296 1492 2304
rect 1644 2296 1652 2304
rect 1724 2296 1732 2304
rect 1836 2296 1844 2304
rect 1884 2296 1892 2304
rect 1900 2296 1908 2304
rect 1980 2296 1988 2304
rect 2156 2296 2164 2304
rect 2188 2296 2196 2304
rect 2348 2296 2356 2304
rect 2412 2296 2420 2304
rect 2476 2296 2484 2304
rect 2556 2296 2564 2304
rect 2620 2296 2628 2304
rect 2652 2296 2660 2304
rect 2700 2296 2708 2304
rect 2764 2296 2772 2304
rect 2844 2296 2852 2304
rect 2908 2296 2916 2304
rect 3164 2316 3172 2324
rect 3228 2316 3236 2324
rect 3260 2316 3268 2324
rect 3292 2316 3300 2324
rect 3388 2316 3396 2324
rect 3468 2316 3476 2324
rect 3532 2316 3540 2324
rect 3580 2316 3588 2324
rect 3660 2316 3668 2324
rect 3788 2316 3796 2324
rect 3900 2316 3908 2324
rect 3964 2316 3972 2324
rect 3004 2296 3012 2304
rect 3084 2296 3092 2304
rect 3180 2296 3188 2304
rect 3196 2296 3204 2304
rect 3244 2296 3252 2304
rect 3308 2296 3316 2304
rect 3500 2296 3508 2304
rect 44 2276 52 2284
rect 108 2276 116 2284
rect 140 2276 148 2284
rect 204 2276 212 2284
rect 236 2276 244 2284
rect 252 2276 260 2284
rect 380 2276 388 2284
rect 444 2276 452 2284
rect 476 2276 484 2284
rect 540 2280 548 2288
rect 3724 2296 3732 2304
rect 3836 2296 3844 2304
rect 3916 2296 3924 2304
rect 4060 2316 4068 2324
rect 4172 2316 4180 2324
rect 4252 2316 4260 2324
rect 4492 2316 4500 2324
rect 4636 2316 4644 2324
rect 4748 2316 4756 2324
rect 5164 2316 5172 2324
rect 5324 2316 5332 2324
rect 5468 2316 5476 2324
rect 5564 2316 5572 2324
rect 5692 2316 5700 2324
rect 5772 2316 5780 2324
rect 5884 2316 5892 2324
rect 6044 2316 6052 2324
rect 6108 2316 6116 2324
rect 4028 2296 4036 2304
rect 4044 2296 4052 2304
rect 4092 2296 4100 2304
rect 4204 2296 4212 2304
rect 4268 2296 4276 2304
rect 4332 2296 4340 2304
rect 4348 2296 4356 2304
rect 4412 2296 4420 2304
rect 4428 2296 4436 2304
rect 4508 2296 4516 2304
rect 4604 2296 4612 2304
rect 4764 2296 4772 2304
rect 4812 2296 4820 2304
rect 5324 2296 5332 2304
rect 5356 2296 5364 2304
rect 5436 2296 5444 2304
rect 5548 2296 5556 2304
rect 5580 2296 5588 2304
rect 5660 2296 5668 2304
rect 5724 2296 5732 2304
rect 5788 2296 5796 2304
rect 5852 2296 5860 2304
rect 5932 2296 5940 2304
rect 6012 2296 6020 2304
rect 6076 2296 6084 2304
rect 556 2276 564 2284
rect 588 2276 596 2284
rect 700 2276 708 2284
rect 796 2276 804 2284
rect 812 2276 820 2284
rect 908 2276 916 2284
rect 1036 2276 1044 2284
rect 1068 2276 1076 2284
rect 1148 2276 1156 2284
rect 1244 2276 1252 2284
rect 1420 2276 1428 2284
rect 1500 2276 1508 2284
rect 1564 2276 1572 2284
rect 1772 2276 1780 2284
rect 1788 2276 1796 2284
rect 1884 2276 1892 2284
rect 2044 2276 2052 2284
rect 2092 2276 2100 2284
rect 2172 2276 2180 2284
rect 2204 2276 2212 2284
rect 2252 2276 2260 2284
rect 2268 2276 2276 2284
rect 2412 2276 2420 2284
rect 2956 2276 2964 2284
rect 2988 2276 2996 2284
rect 3068 2276 3076 2284
rect 3132 2276 3140 2284
rect 3244 2276 3252 2284
rect 3356 2276 3364 2284
rect 3436 2276 3444 2284
rect 3484 2276 3492 2284
rect 3516 2276 3524 2284
rect 3564 2276 3572 2284
rect 3612 2276 3620 2284
rect 3628 2276 3636 2284
rect 3964 2276 3972 2284
rect 4012 2276 4020 2284
rect 4076 2276 4084 2284
rect 4140 2276 4148 2284
rect 4188 2276 4196 2284
rect 4364 2276 4372 2284
rect 4396 2276 4404 2284
rect 156 2256 164 2264
rect 412 2256 420 2264
rect 620 2256 628 2264
rect 876 2256 884 2264
rect 940 2256 948 2264
rect 1308 2256 1316 2264
rect 1388 2256 1396 2264
rect 1804 2256 1812 2264
rect 2108 2256 2116 2264
rect 2252 2256 2260 2264
rect 2508 2256 2516 2264
rect 2812 2256 2820 2264
rect 3052 2256 3060 2264
rect 3276 2256 3284 2264
rect 3452 2256 3460 2264
rect 3724 2256 3732 2264
rect 3884 2256 3892 2264
rect 4316 2256 4324 2264
rect 4460 2256 4468 2264
rect 4540 2256 4548 2264
rect 4572 2276 4580 2284
rect 4588 2276 4596 2284
rect 4652 2276 4660 2284
rect 4700 2276 4708 2284
rect 4764 2276 4772 2284
rect 4828 2276 4836 2284
rect 4940 2276 4948 2284
rect 4988 2280 4996 2288
rect 5004 2276 5012 2284
rect 5020 2276 5028 2284
rect 5052 2276 5060 2284
rect 5116 2276 5124 2284
rect 5180 2276 5188 2284
rect 5276 2276 5284 2284
rect 5292 2276 5300 2284
rect 5324 2276 5332 2284
rect 5468 2276 5476 2284
rect 5500 2276 5508 2284
rect 5596 2276 5604 2284
rect 5644 2276 5652 2284
rect 5708 2276 5716 2284
rect 6060 2276 6068 2284
rect 6124 2276 6132 2284
rect 6236 2276 6244 2284
rect 5116 2256 5124 2264
rect 5148 2256 5156 2264
rect 5468 2256 5476 2264
rect 5628 2256 5636 2264
rect 5932 2256 5940 2264
rect 5980 2256 5988 2264
rect 28 2236 36 2244
rect 76 2236 84 2244
rect 108 2236 116 2244
rect 332 2236 340 2244
rect 396 2236 404 2244
rect 476 2236 484 2244
rect 508 2236 516 2244
rect 748 2236 756 2244
rect 764 2236 772 2244
rect 860 2236 868 2244
rect 956 2236 964 2244
rect 1180 2236 1188 2244
rect 1260 2236 1268 2244
rect 1356 2236 1364 2244
rect 1404 2236 1412 2244
rect 1516 2236 1524 2244
rect 1676 2236 1684 2244
rect 1724 2236 1732 2244
rect 2028 2236 2036 2244
rect 2060 2236 2068 2244
rect 2300 2236 2308 2244
rect 2876 2236 2884 2244
rect 2988 2236 2996 2244
rect 3036 2236 3044 2244
rect 3388 2236 3396 2244
rect 3548 2236 3556 2244
rect 4172 2236 4180 2244
rect 4236 2236 4244 2244
rect 4268 2236 4276 2244
rect 4396 2236 4404 2244
rect 4748 2236 4756 2244
rect 4908 2236 4916 2244
rect 4956 2236 4964 2244
rect 5052 2236 5060 2244
rect 5068 2236 5076 2244
rect 5756 2236 5764 2244
rect 5852 2236 5860 2244
rect 6156 2236 6164 2244
rect 3118 2206 3126 2214
rect 3132 2206 3140 2214
rect 3146 2206 3154 2214
rect 508 2176 516 2184
rect 684 2176 692 2184
rect 956 2176 964 2184
rect 1196 2176 1204 2184
rect 1948 2176 1956 2184
rect 2412 2176 2420 2184
rect 2668 2176 2676 2184
rect 2748 2176 2756 2184
rect 2956 2176 2964 2184
rect 2988 2176 2996 2184
rect 3036 2176 3044 2184
rect 3292 2176 3300 2184
rect 3516 2176 3524 2184
rect 3852 2176 3860 2184
rect 4236 2176 4244 2184
rect 4444 2176 4452 2184
rect 4508 2176 4516 2184
rect 4684 2176 4692 2184
rect 4780 2176 4788 2184
rect 5132 2176 5140 2184
rect 5212 2176 5220 2184
rect 5788 2176 5796 2184
rect 5868 2176 5876 2184
rect 6012 2176 6020 2184
rect 6236 2176 6244 2184
rect 156 2156 164 2164
rect 172 2156 180 2164
rect 300 2156 308 2164
rect 748 2156 756 2164
rect 908 2156 916 2164
rect 1212 2156 1220 2164
rect 1228 2156 1236 2164
rect 1276 2156 1284 2164
rect 1756 2156 1764 2164
rect 1964 2156 1972 2164
rect 2092 2156 2100 2164
rect 2396 2156 2404 2164
rect 2572 2156 2580 2164
rect 2892 2156 2900 2164
rect 3052 2156 3060 2164
rect 3372 2156 3380 2164
rect 3532 2156 3540 2164
rect 3564 2156 3572 2164
rect 3580 2156 3588 2164
rect 172 2136 180 2144
rect 204 2132 212 2140
rect 268 2136 276 2144
rect 380 2136 388 2144
rect 556 2136 564 2144
rect 716 2136 724 2144
rect 844 2136 852 2144
rect 876 2136 884 2144
rect 972 2136 980 2144
rect 1068 2136 1076 2144
rect 1404 2136 1412 2144
rect 1436 2136 1444 2144
rect 1916 2136 1924 2144
rect 1996 2136 2004 2144
rect 2124 2136 2132 2144
rect 2364 2136 2372 2144
rect 2508 2136 2516 2144
rect 2524 2136 2532 2144
rect 2572 2136 2580 2144
rect 2604 2136 2612 2144
rect 2684 2136 2692 2144
rect 2796 2136 2804 2144
rect 2812 2136 2820 2144
rect 2844 2136 2852 2144
rect 3004 2136 3012 2144
rect 3244 2136 3252 2144
rect 3308 2136 3316 2144
rect 3404 2136 3412 2144
rect 3436 2136 3444 2144
rect 3452 2136 3460 2144
rect 3468 2132 3476 2140
rect 3596 2136 3604 2144
rect 3708 2136 3716 2144
rect 3740 2136 3748 2144
rect 3868 2156 3876 2164
rect 4012 2156 4020 2164
rect 4220 2156 4228 2164
rect 4732 2156 4740 2164
rect 3900 2136 3908 2144
rect 3948 2136 3956 2144
rect 3964 2136 3972 2144
rect 4028 2136 4036 2144
rect 4252 2136 4260 2144
rect 4284 2136 4292 2144
rect 4348 2136 4356 2144
rect 4396 2136 4404 2144
rect 4460 2136 4468 2144
rect 5068 2156 5076 2164
rect 5164 2156 5172 2164
rect 5628 2156 5636 2164
rect 6252 2156 6260 2164
rect 4828 2136 4836 2144
rect 4844 2136 4852 2144
rect 4940 2136 4948 2144
rect 5036 2136 5044 2144
rect 5100 2136 5108 2144
rect 5148 2136 5156 2144
rect 5228 2136 5236 2144
rect 5324 2136 5332 2144
rect 5388 2136 5396 2144
rect 5580 2136 5588 2144
rect 5628 2136 5636 2144
rect 5660 2136 5668 2144
rect 5772 2136 5780 2144
rect 5836 2136 5844 2144
rect 5884 2136 5892 2144
rect 6028 2136 6036 2144
rect 6124 2136 6132 2144
rect 6140 2136 6148 2144
rect 6204 2136 6212 2144
rect 6220 2136 6228 2144
rect 44 2116 52 2124
rect 92 2116 100 2124
rect 140 2116 148 2124
rect 236 2116 244 2124
rect 252 2116 260 2124
rect 316 2116 324 2124
rect 380 2116 388 2124
rect 428 2116 436 2124
rect 476 2116 484 2124
rect 540 2116 548 2124
rect 604 2116 612 2124
rect 652 2116 660 2124
rect 700 2116 708 2124
rect 780 2116 788 2124
rect 828 2116 836 2124
rect 908 2116 916 2124
rect 988 2116 996 2124
rect 1020 2116 1028 2124
rect 1180 2116 1188 2124
rect 1308 2116 1316 2124
rect 1356 2116 1364 2124
rect 1420 2116 1428 2124
rect 1500 2116 1508 2124
rect 1532 2116 1540 2124
rect 1644 2116 1652 2124
rect 1724 2116 1732 2124
rect 1804 2116 1812 2124
rect 1868 2116 1876 2124
rect 2012 2116 2020 2124
rect 2044 2116 2052 2124
rect 2140 2116 2148 2124
rect 2172 2116 2180 2124
rect 2204 2116 2212 2124
rect 2252 2116 2260 2124
rect 2300 2116 2308 2124
rect 2348 2116 2356 2124
rect 2412 2116 2420 2124
rect 2444 2116 2452 2124
rect 60 2096 68 2104
rect 76 2096 84 2104
rect 364 2096 372 2104
rect 428 2096 436 2104
rect 492 2096 500 2104
rect 508 2096 516 2104
rect 620 2096 628 2104
rect 636 2096 644 2104
rect 780 2096 788 2104
rect 1004 2096 1012 2104
rect 1372 2096 1380 2104
rect 1388 2096 1396 2104
rect 1500 2096 1508 2104
rect 1516 2096 1524 2104
rect 1628 2096 1636 2104
rect 1852 2096 1860 2104
rect 1900 2096 1908 2104
rect 1948 2096 1956 2104
rect 2028 2096 2036 2104
rect 2076 2096 2084 2104
rect 2156 2096 2164 2104
rect 2268 2096 2276 2104
rect 2412 2096 2420 2104
rect 2476 2096 2484 2104
rect 2556 2096 2564 2104
rect 2636 2096 2644 2104
rect 2780 2116 2788 2124
rect 2924 2116 2932 2124
rect 3004 2116 3012 2124
rect 3100 2116 3108 2124
rect 3196 2116 3204 2124
rect 3260 2116 3268 2124
rect 3420 2116 3428 2124
rect 3676 2116 3684 2124
rect 3772 2116 3780 2124
rect 3788 2116 3796 2124
rect 3820 2116 3828 2124
rect 3900 2116 3908 2124
rect 3916 2116 3924 2124
rect 3980 2116 3988 2124
rect 4044 2116 4052 2124
rect 4076 2116 4084 2124
rect 4108 2116 4116 2124
rect 4188 2116 4196 2124
rect 4268 2116 4276 2124
rect 4300 2116 4308 2124
rect 4396 2116 4404 2124
rect 4412 2116 4420 2124
rect 4476 2116 4484 2124
rect 4540 2116 4548 2124
rect 4604 2116 4612 2124
rect 4668 2116 4676 2124
rect 4700 2116 4708 2124
rect 4812 2116 4820 2124
rect 4940 2116 4948 2124
rect 4972 2116 4980 2124
rect 5020 2116 5028 2124
rect 5068 2116 5076 2124
rect 5084 2116 5092 2124
rect 5148 2116 5156 2124
rect 5244 2116 5252 2124
rect 5292 2116 5300 2124
rect 5340 2116 5348 2124
rect 5388 2116 5396 2124
rect 5404 2116 5412 2124
rect 5420 2116 5428 2124
rect 5484 2116 5492 2124
rect 5532 2116 5540 2124
rect 5564 2116 5572 2124
rect 5676 2116 5684 2124
rect 5724 2116 5732 2124
rect 5980 2116 5988 2124
rect 6044 2116 6052 2124
rect 6076 2116 6084 2124
rect 6124 2116 6132 2124
rect 6188 2116 6196 2124
rect 6204 2116 6212 2124
rect 2732 2096 2740 2104
rect 2892 2096 2900 2104
rect 2908 2096 2916 2104
rect 2972 2096 2980 2104
rect 3068 2096 3076 2104
rect 3228 2096 3236 2104
rect 3340 2096 3348 2104
rect 3356 2096 3364 2104
rect 3388 2096 3396 2104
rect 3676 2096 3684 2104
rect 3708 2096 3716 2104
rect 3948 2096 3956 2104
rect 4012 2096 4020 2104
rect 4140 2096 4148 2104
rect 4204 2096 4212 2104
rect 4380 2096 4388 2104
rect 4444 2096 4452 2104
rect 4508 2096 4516 2104
rect 4524 2096 4532 2104
rect 4588 2096 4596 2104
rect 4860 2096 4868 2104
rect 4876 2096 4884 2104
rect 4892 2096 4900 2104
rect 5004 2096 5012 2104
rect 5308 2096 5316 2104
rect 5372 2096 5380 2104
rect 5436 2096 5444 2104
rect 5500 2096 5508 2104
rect 5516 2096 5524 2104
rect 5612 2096 5620 2104
rect 5740 2096 5748 2104
rect 5884 2096 5892 2104
rect 5932 2096 5940 2104
rect 6060 2096 6068 2104
rect 6172 2096 6180 2104
rect 28 2076 36 2084
rect 108 2076 116 2084
rect 460 2076 468 2084
rect 764 2076 772 2084
rect 1036 2076 1044 2084
rect 1260 2076 1268 2084
rect 1308 2076 1316 2084
rect 1324 2076 1332 2084
rect 1340 2076 1348 2084
rect 1356 2076 1364 2084
rect 1644 2076 1652 2084
rect 1660 2076 1668 2084
rect 1708 2076 1716 2084
rect 1820 2076 1828 2084
rect 1884 2076 1892 2084
rect 2060 2076 2068 2084
rect 2188 2076 2196 2084
rect 2236 2076 2244 2084
rect 2252 2076 2260 2084
rect 2572 2076 2580 2084
rect 2812 2076 2820 2084
rect 2924 2076 2932 2084
rect 2940 2076 2948 2084
rect 3084 2076 3092 2084
rect 3196 2076 3204 2084
rect 300 2056 308 2064
rect 476 2056 484 2064
rect 1100 2056 1108 2064
rect 3244 2076 3252 2084
rect 3500 2076 3508 2084
rect 3564 2076 3572 2084
rect 3628 2076 3636 2084
rect 3660 2076 3668 2084
rect 4108 2076 4116 2084
rect 4172 2076 4180 2084
rect 4348 2076 4356 2084
rect 4556 2076 4564 2084
rect 4604 2076 4612 2084
rect 4620 2076 4628 2084
rect 4988 2076 4996 2084
rect 5276 2076 5284 2084
rect 5468 2076 5476 2084
rect 5484 2076 5492 2084
rect 5708 2076 5716 2084
rect 6092 2076 6100 2084
rect 4188 2056 4196 2064
rect 5292 2056 5300 2064
rect 5724 2056 5732 2064
rect 12 2036 20 2044
rect 124 2036 132 2044
rect 332 2036 340 2044
rect 748 2036 756 2044
rect 812 2036 820 2044
rect 876 2036 884 2044
rect 1052 2036 1060 2044
rect 1676 2036 1684 2044
rect 1724 2036 1732 2044
rect 1804 2036 1812 2044
rect 1868 2036 1876 2044
rect 1964 2036 1972 2044
rect 2092 2036 2100 2044
rect 2220 2036 2228 2044
rect 2332 2036 2340 2044
rect 2492 2036 2500 2044
rect 2716 2036 2724 2044
rect 3164 2036 3172 2044
rect 3324 2036 3332 2044
rect 3676 2036 3684 2044
rect 4092 2036 4100 2044
rect 4764 2036 4772 2044
rect 4924 2036 4932 2044
rect 4988 2036 4996 2044
rect 5452 2036 5460 2044
rect 5596 2036 5604 2044
rect 5628 2036 5636 2044
rect 1566 2006 1574 2014
rect 1580 2006 1588 2014
rect 1594 2006 1602 2014
rect 4638 2006 4646 2014
rect 4652 2006 4660 2014
rect 4666 2006 4674 2014
rect 460 1976 468 1984
rect 828 1976 836 1984
rect 908 1976 916 1984
rect 972 1976 980 1984
rect 1116 1976 1124 1984
rect 1292 1976 1300 1984
rect 1420 1976 1428 1984
rect 1756 1976 1764 1984
rect 2380 1976 2388 1984
rect 2444 1976 2452 1984
rect 2524 1976 2532 1984
rect 2588 1976 2596 1984
rect 2620 1976 2628 1984
rect 3276 1976 3284 1984
rect 3436 1976 3444 1984
rect 3628 1976 3636 1984
rect 3916 1976 3924 1984
rect 5772 1976 5780 1984
rect 6220 1976 6228 1984
rect 1372 1956 1380 1964
rect 2060 1956 2068 1964
rect 2972 1956 2980 1964
rect 268 1936 276 1944
rect 300 1936 308 1944
rect 1100 1936 1108 1944
rect 1228 1936 1236 1944
rect 1260 1936 1268 1944
rect 1356 1936 1364 1944
rect 1772 1936 1780 1944
rect 2044 1936 2052 1944
rect 2172 1936 2180 1944
rect 2364 1936 2372 1944
rect 2476 1936 2484 1944
rect 2508 1936 2516 1944
rect 2636 1936 2644 1944
rect 2716 1936 2724 1944
rect 2764 1936 2772 1944
rect 2796 1936 2804 1944
rect 2956 1936 2964 1944
rect 2988 1936 2996 1944
rect 3084 1936 3092 1944
rect 4412 1956 4420 1964
rect 5484 1956 5492 1964
rect 5948 1956 5956 1964
rect 3148 1936 3156 1944
rect 3164 1936 3172 1944
rect 3260 1936 3268 1944
rect 3324 1936 3332 1944
rect 3932 1936 3940 1944
rect 4316 1936 4324 1944
rect 4444 1936 4452 1944
rect 4780 1936 4788 1944
rect 4812 1936 4820 1944
rect 5468 1936 5476 1944
rect 5692 1936 5700 1944
rect 5756 1936 5764 1944
rect 5852 1936 5860 1944
rect 5932 1936 5940 1944
rect 5996 1936 6004 1944
rect 332 1916 340 1924
rect 476 1916 484 1924
rect 12 1896 20 1904
rect 76 1896 84 1904
rect 140 1896 148 1904
rect 156 1896 164 1904
rect 220 1896 228 1904
rect 284 1896 292 1904
rect 396 1896 404 1904
rect 476 1896 484 1904
rect 588 1916 596 1924
rect 636 1916 644 1924
rect 668 1916 676 1924
rect 796 1916 804 1924
rect 812 1916 820 1924
rect 1004 1916 1012 1924
rect 1068 1916 1076 1924
rect 1132 1916 1140 1924
rect 1212 1916 1220 1924
rect 1324 1916 1332 1924
rect 1388 1916 1396 1924
rect 1644 1916 1652 1924
rect 1724 1916 1732 1924
rect 1740 1916 1748 1924
rect 1868 1916 1876 1924
rect 1900 1916 1908 1924
rect 1932 1916 1940 1924
rect 2012 1916 2020 1924
rect 2076 1916 2084 1924
rect 2204 1916 2212 1924
rect 2396 1916 2404 1924
rect 2460 1916 2468 1924
rect 2604 1916 2612 1924
rect 2716 1916 2724 1924
rect 2732 1916 2740 1924
rect 2844 1916 2852 1924
rect 2892 1916 2900 1924
rect 2924 1916 2932 1924
rect 2988 1916 2996 1924
rect 3116 1916 3124 1924
rect 3292 1916 3300 1924
rect 3516 1916 3524 1924
rect 3676 1916 3684 1924
rect 3708 1916 3716 1924
rect 3740 1916 3748 1924
rect 3820 1916 3828 1924
rect 3868 1916 3876 1924
rect 3932 1916 3940 1924
rect 4012 1916 4020 1924
rect 4188 1916 4196 1924
rect 4284 1916 4292 1924
rect 4348 1916 4356 1924
rect 4364 1916 4372 1924
rect 4476 1916 4484 1924
rect 4556 1916 4564 1924
rect 4844 1916 4852 1924
rect 4924 1916 4932 1924
rect 5180 1916 5188 1924
rect 5196 1916 5204 1924
rect 684 1896 692 1904
rect 748 1896 756 1904
rect 876 1896 884 1904
rect 940 1896 948 1904
rect 1004 1896 1012 1904
rect 1116 1896 1124 1904
rect 1148 1896 1156 1904
rect 1196 1896 1204 1904
rect 1228 1896 1236 1904
rect 1292 1896 1300 1904
rect 1372 1896 1380 1904
rect 1436 1896 1444 1904
rect 1500 1896 1508 1904
rect 1516 1896 1524 1904
rect 1756 1896 1764 1904
rect 1804 1896 1812 1904
rect 1964 1896 1972 1904
rect 2012 1896 2020 1904
rect 2060 1896 2068 1904
rect 2092 1896 2100 1904
rect 2188 1896 2196 1904
rect 2220 1896 2228 1904
rect 2316 1896 2324 1904
rect 2380 1896 2388 1904
rect 2444 1896 2452 1904
rect 2492 1896 2500 1904
rect 2540 1896 2548 1904
rect 2620 1896 2628 1904
rect 2700 1896 2708 1904
rect 2748 1896 2756 1904
rect 2972 1896 2980 1904
rect 3004 1896 3012 1904
rect 3100 1896 3108 1904
rect 3164 1896 3172 1904
rect 3276 1896 3284 1904
rect 3340 1896 3348 1904
rect 3436 1896 3444 1904
rect 3628 1896 3636 1904
rect 3644 1896 3652 1904
rect 3724 1896 3732 1904
rect 3916 1896 3924 1904
rect 3948 1896 3956 1904
rect 4060 1896 4068 1904
rect 4124 1896 4132 1904
rect 4156 1896 4164 1904
rect 4204 1896 4212 1904
rect 4220 1896 4228 1904
rect 4332 1896 4340 1904
rect 4380 1896 4388 1904
rect 4460 1896 4468 1904
rect 4492 1896 4500 1904
rect 4604 1896 4612 1904
rect 28 1876 36 1884
rect 92 1876 100 1884
rect 172 1876 180 1884
rect 204 1876 212 1884
rect 364 1876 372 1884
rect 380 1876 388 1884
rect 444 1876 452 1884
rect 524 1876 532 1884
rect 572 1876 580 1884
rect 636 1876 644 1884
rect 684 1876 692 1884
rect 732 1876 740 1884
rect 764 1876 772 1884
rect 860 1876 868 1884
rect 956 1876 964 1884
rect 1020 1876 1028 1884
rect 1164 1876 1172 1884
rect 1276 1876 1284 1884
rect 1452 1876 1460 1884
rect 1484 1876 1492 1884
rect 1516 1876 1524 1884
rect 1564 1876 1572 1884
rect 1676 1876 1684 1884
rect 1692 1876 1700 1884
rect 1724 1876 1732 1884
rect 1820 1876 1828 1884
rect 60 1856 68 1864
rect 236 1856 244 1864
rect 940 1856 948 1864
rect 1196 1856 1204 1864
rect 1404 1856 1412 1864
rect 1644 1856 1652 1864
rect 1948 1876 1956 1884
rect 2108 1876 2116 1884
rect 2236 1876 2244 1884
rect 2332 1876 2340 1884
rect 2556 1876 2564 1884
rect 2684 1876 2692 1884
rect 2844 1876 2852 1884
rect 2892 1876 2900 1884
rect 3020 1876 3028 1884
rect 3196 1876 3204 1884
rect 3452 1876 3460 1884
rect 3548 1876 3556 1884
rect 3644 1876 3652 1884
rect 3660 1876 3668 1884
rect 3724 1876 3732 1884
rect 3788 1876 3796 1884
rect 3836 1876 3844 1884
rect 3964 1876 3972 1884
rect 4828 1896 4836 1904
rect 4876 1896 4884 1904
rect 4924 1896 4932 1904
rect 4956 1896 4964 1904
rect 5020 1896 5028 1904
rect 4076 1876 4084 1884
rect 4108 1876 4116 1884
rect 4124 1876 4132 1884
rect 4204 1876 4212 1884
rect 4252 1876 4260 1884
rect 4508 1876 4516 1884
rect 4588 1876 4596 1884
rect 4620 1876 4628 1884
rect 4652 1876 4660 1884
rect 4732 1876 4740 1884
rect 4748 1880 4756 1888
rect 4860 1876 4868 1884
rect 4940 1876 4948 1884
rect 5036 1876 5044 1884
rect 5148 1896 5156 1904
rect 5324 1896 5332 1904
rect 5548 1916 5556 1924
rect 5580 1916 5588 1924
rect 5660 1916 5668 1924
rect 5724 1916 5732 1924
rect 5788 1916 5796 1924
rect 5884 1916 5892 1924
rect 5900 1916 5908 1924
rect 5964 1916 5972 1924
rect 6028 1916 6036 1924
rect 5372 1896 5380 1904
rect 5436 1896 5444 1904
rect 5484 1896 5492 1904
rect 5628 1896 5636 1904
rect 5708 1896 5716 1904
rect 5772 1896 5780 1904
rect 5868 1896 5876 1904
rect 5916 1896 5924 1904
rect 5980 1896 5988 1904
rect 6108 1896 6116 1904
rect 6172 1896 6180 1904
rect 6236 1896 6244 1904
rect 5148 1876 5156 1884
rect 5228 1876 5236 1884
rect 5244 1876 5252 1884
rect 5276 1876 5284 1884
rect 5388 1876 5396 1884
rect 5420 1876 5428 1884
rect 5596 1876 5604 1884
rect 5660 1876 5668 1884
rect 5708 1876 5716 1884
rect 5868 1876 5876 1884
rect 6028 1876 6036 1884
rect 6060 1876 6068 1884
rect 6092 1876 6100 1884
rect 6188 1876 6196 1884
rect 6236 1876 6244 1884
rect 1868 1856 1876 1864
rect 2140 1856 2148 1864
rect 2268 1856 2276 1864
rect 2588 1856 2596 1864
rect 3036 1856 3044 1864
rect 3052 1856 3060 1864
rect 3228 1856 3236 1864
rect 3388 1856 3396 1864
rect 3532 1856 3540 1864
rect 3980 1856 3988 1864
rect 3996 1856 4004 1864
rect 4108 1856 4116 1864
rect 4284 1856 4292 1864
rect 4332 1856 4340 1864
rect 4540 1856 4548 1864
rect 4828 1856 4836 1864
rect 4988 1856 4996 1864
rect 5180 1856 5188 1864
rect 5292 1856 5300 1864
rect 5356 1856 5364 1864
rect 5420 1856 5428 1864
rect 5532 1856 5540 1864
rect 5804 1856 5812 1864
rect 6156 1856 6164 1864
rect 44 1836 52 1844
rect 124 1836 132 1844
rect 188 1836 196 1844
rect 284 1836 292 1844
rect 348 1836 356 1844
rect 492 1836 500 1844
rect 508 1836 516 1844
rect 572 1836 580 1844
rect 620 1836 628 1844
rect 668 1836 676 1844
rect 716 1836 724 1844
rect 780 1836 788 1844
rect 812 1836 820 1844
rect 908 1836 916 1844
rect 924 1836 932 1844
rect 1068 1836 1076 1844
rect 1468 1836 1476 1844
rect 1532 1836 1540 1844
rect 2124 1836 2132 1844
rect 2172 1836 2180 1844
rect 2252 1836 2260 1844
rect 2284 1836 2292 1844
rect 2812 1836 2820 1844
rect 2924 1836 2932 1844
rect 3212 1836 3220 1844
rect 3340 1836 3348 1844
rect 3516 1836 3524 1844
rect 3820 1836 3828 1844
rect 3868 1836 3876 1844
rect 4460 1836 4468 1844
rect 4524 1836 4532 1844
rect 4620 1836 4628 1844
rect 5068 1836 5076 1844
rect 5196 1836 5204 1844
rect 5820 1836 5828 1844
rect 6028 1836 6036 1844
rect 3118 1806 3126 1814
rect 3132 1806 3140 1814
rect 3146 1806 3154 1814
rect 92 1776 100 1784
rect 140 1776 148 1784
rect 396 1776 404 1784
rect 2156 1776 2164 1784
rect 2364 1776 2372 1784
rect 2444 1776 2452 1784
rect 2556 1776 2564 1784
rect 2812 1776 2820 1784
rect 2892 1776 2900 1784
rect 2972 1776 2980 1784
rect 3308 1776 3316 1784
rect 3436 1776 3444 1784
rect 3708 1776 3716 1784
rect 4572 1776 4580 1784
rect 4812 1776 4820 1784
rect 4876 1776 4884 1784
rect 5132 1776 5140 1784
rect 5212 1776 5220 1784
rect 5276 1776 5284 1784
rect 5340 1776 5348 1784
rect 5548 1776 5556 1784
rect 5788 1776 5796 1784
rect 6252 1776 6260 1784
rect 300 1756 308 1764
rect 380 1756 388 1764
rect 524 1756 532 1764
rect 796 1756 804 1764
rect 1068 1756 1076 1764
rect 1196 1756 1204 1764
rect 1420 1756 1428 1764
rect 1996 1756 2004 1764
rect 2524 1756 2532 1764
rect 2796 1756 2804 1764
rect 2908 1756 2916 1764
rect 3004 1756 3012 1764
rect 3100 1756 3108 1764
rect 3212 1756 3220 1764
rect 3276 1756 3284 1764
rect 3292 1756 3300 1764
rect 3388 1756 3396 1764
rect 3500 1756 3508 1764
rect 3564 1756 3572 1764
rect 3628 1756 3636 1764
rect 3932 1756 3940 1764
rect 4012 1756 4020 1764
rect 4076 1756 4084 1764
rect 444 1736 452 1744
rect 460 1736 468 1744
rect 476 1732 484 1740
rect 556 1736 564 1744
rect 636 1736 644 1744
rect 684 1736 692 1744
rect 716 1736 724 1744
rect 748 1736 756 1744
rect 796 1736 804 1744
rect 892 1736 900 1744
rect 940 1736 948 1744
rect 988 1736 996 1744
rect 1020 1736 1028 1744
rect 1052 1736 1060 1744
rect 1100 1736 1108 1744
rect 1116 1736 1124 1744
rect 1148 1736 1156 1744
rect 1244 1736 1252 1744
rect 1308 1736 1316 1744
rect 1372 1736 1380 1744
rect 1436 1736 1444 1744
rect 1484 1736 1492 1744
rect 1596 1736 1604 1744
rect 1660 1736 1668 1744
rect 1708 1736 1716 1744
rect 1724 1736 1732 1744
rect 1772 1736 1780 1744
rect 1884 1736 1892 1744
rect 2060 1736 2068 1744
rect 2252 1736 2260 1744
rect 2620 1736 2628 1744
rect 2748 1736 2756 1744
rect 2812 1736 2820 1744
rect 2844 1736 2852 1744
rect 2908 1736 2916 1744
rect 3180 1736 3188 1744
rect 3260 1736 3268 1744
rect 3356 1736 3364 1744
rect 3612 1736 3620 1744
rect 3692 1736 3700 1744
rect 3740 1736 3748 1744
rect 12 1716 20 1724
rect 60 1716 68 1724
rect 108 1716 116 1724
rect 156 1716 164 1724
rect 236 1716 244 1724
rect 268 1716 276 1724
rect 332 1716 340 1724
rect 412 1716 420 1724
rect 508 1716 516 1724
rect 556 1716 564 1724
rect 668 1716 676 1724
rect 700 1716 708 1724
rect 732 1716 740 1724
rect 844 1716 852 1724
rect 876 1716 884 1724
rect 940 1716 948 1724
rect 1036 1716 1044 1724
rect 1244 1716 1252 1724
rect 1292 1716 1300 1724
rect 1356 1716 1364 1724
rect 1388 1716 1396 1724
rect 1420 1716 1428 1724
rect 1468 1716 1476 1724
rect 1532 1716 1540 1724
rect 1644 1716 1652 1724
rect 1788 1716 1796 1724
rect 252 1696 260 1704
rect 332 1696 340 1704
rect 412 1696 420 1704
rect 588 1696 596 1704
rect 764 1696 772 1704
rect 956 1696 964 1704
rect 1004 1696 1012 1704
rect 1132 1696 1140 1704
rect 1196 1696 1204 1704
rect 1260 1696 1268 1704
rect 1468 1696 1476 1704
rect 1548 1696 1556 1704
rect 1676 1696 1684 1704
rect 1756 1696 1764 1704
rect 1868 1716 1876 1724
rect 1932 1716 1940 1724
rect 1964 1716 1972 1724
rect 2044 1716 2052 1724
rect 2108 1716 2116 1724
rect 2172 1716 2180 1724
rect 2220 1716 2228 1724
rect 2236 1716 2244 1724
rect 2364 1716 2372 1724
rect 2412 1716 2420 1724
rect 2476 1716 2484 1724
rect 2588 1716 2596 1724
rect 2636 1716 2644 1724
rect 2668 1716 2676 1724
rect 2716 1716 2724 1724
rect 2748 1716 2756 1724
rect 2860 1716 2868 1724
rect 2940 1716 2948 1724
rect 2972 1716 2980 1724
rect 3052 1716 3060 1724
rect 3100 1716 3108 1724
rect 3228 1716 3236 1724
rect 3340 1716 3348 1724
rect 3548 1716 3556 1724
rect 3676 1716 3684 1724
rect 3740 1716 3748 1724
rect 3868 1736 3876 1744
rect 4060 1736 4068 1744
rect 4140 1736 4148 1744
rect 4188 1736 4196 1744
rect 4204 1736 4212 1744
rect 4316 1736 4324 1744
rect 4364 1736 4372 1744
rect 4476 1736 4484 1744
rect 4588 1756 4596 1764
rect 4732 1756 4740 1764
rect 4924 1756 4932 1764
rect 4604 1736 4612 1744
rect 4796 1736 4804 1744
rect 4828 1736 4836 1744
rect 5356 1756 5364 1764
rect 5564 1756 5572 1764
rect 5596 1756 5604 1764
rect 5708 1756 5716 1764
rect 4972 1736 4980 1744
rect 5068 1736 5076 1744
rect 5084 1736 5092 1744
rect 5148 1736 5156 1744
rect 5260 1736 5268 1744
rect 5292 1736 5300 1744
rect 5308 1736 5316 1744
rect 5500 1736 5508 1744
rect 5516 1732 5524 1740
rect 5628 1736 5636 1744
rect 5724 1736 5732 1744
rect 3772 1716 3780 1724
rect 1836 1696 1844 1704
rect 1868 1696 1876 1704
rect 252 1676 260 1684
rect 348 1676 356 1684
rect 828 1676 836 1684
rect 1164 1676 1172 1684
rect 1916 1676 1924 1684
rect 2012 1696 2020 1704
rect 2124 1696 2132 1704
rect 2188 1696 2196 1704
rect 2204 1696 2212 1704
rect 2316 1696 2324 1704
rect 2380 1696 2388 1704
rect 2092 1676 2100 1684
rect 2156 1676 2164 1684
rect 2284 1676 2292 1684
rect 2348 1676 2356 1684
rect 2364 1676 2372 1684
rect 2460 1696 2468 1704
rect 2604 1696 2612 1704
rect 2668 1696 2676 1704
rect 2732 1696 2740 1704
rect 2812 1696 2820 1704
rect 2972 1696 2980 1704
rect 3068 1696 3076 1704
rect 3228 1696 3236 1704
rect 3644 1696 3652 1704
rect 3708 1696 3716 1704
rect 3804 1696 3812 1704
rect 3852 1716 3860 1724
rect 3980 1716 3988 1724
rect 4124 1716 4132 1724
rect 4140 1716 4148 1724
rect 4220 1716 4228 1724
rect 4236 1716 4244 1724
rect 4092 1696 4100 1704
rect 4156 1696 4164 1704
rect 4300 1716 4308 1724
rect 4268 1696 4276 1704
rect 4332 1696 4340 1704
rect 4412 1696 4420 1704
rect 4476 1716 4484 1724
rect 4524 1716 4532 1724
rect 4588 1716 4596 1724
rect 4700 1716 4708 1724
rect 4732 1716 4740 1724
rect 4764 1716 4772 1724
rect 4892 1716 4900 1724
rect 4988 1716 4996 1724
rect 4748 1696 4756 1704
rect 4876 1696 4884 1704
rect 4908 1696 4916 1704
rect 5308 1716 5316 1724
rect 5388 1716 5396 1724
rect 5420 1716 5428 1724
rect 5468 1716 5476 1724
rect 5644 1716 5652 1724
rect 5708 1716 5716 1724
rect 5740 1716 5748 1724
rect 5916 1736 5924 1744
rect 5948 1736 5956 1744
rect 6172 1736 6180 1744
rect 5852 1716 5860 1724
rect 5980 1718 5988 1726
rect 6044 1716 6052 1724
rect 6124 1716 6132 1724
rect 6188 1716 6196 1724
rect 5036 1696 5044 1704
rect 5132 1696 5140 1704
rect 5260 1696 5268 1704
rect 5372 1696 5380 1704
rect 5484 1696 5492 1704
rect 5596 1696 5604 1704
rect 5676 1696 5684 1704
rect 5884 1696 5892 1704
rect 6236 1696 6244 1704
rect 2428 1676 2436 1684
rect 2460 1676 2468 1684
rect 2540 1676 2548 1684
rect 2572 1676 2580 1684
rect 2700 1676 2708 1684
rect 3036 1676 3044 1684
rect 3052 1676 3060 1684
rect 4348 1676 4356 1684
rect 4780 1676 4788 1684
rect 5404 1676 5412 1684
rect 5452 1676 5460 1684
rect 6108 1676 6116 1684
rect 6156 1676 6164 1684
rect 92 1656 100 1664
rect 1148 1656 1156 1664
rect 1324 1656 1332 1664
rect 1612 1656 1620 1664
rect 1692 1656 1700 1664
rect 2108 1656 2116 1664
rect 4028 1656 4036 1664
rect 4396 1656 4404 1664
rect 4956 1656 4964 1664
rect 44 1636 52 1644
rect 188 1636 196 1644
rect 236 1636 244 1644
rect 268 1636 276 1644
rect 332 1636 340 1644
rect 572 1636 580 1644
rect 860 1636 868 1644
rect 924 1636 932 1644
rect 1068 1636 1076 1644
rect 1292 1636 1300 1644
rect 1404 1636 1412 1644
rect 1500 1636 1508 1644
rect 1788 1636 1796 1644
rect 1900 1636 1908 1644
rect 2044 1636 2052 1644
rect 2476 1636 2484 1644
rect 2716 1636 2724 1644
rect 2828 1636 2836 1644
rect 3020 1636 3028 1644
rect 3580 1636 3588 1644
rect 3676 1636 3684 1644
rect 3852 1636 3860 1644
rect 3884 1636 3892 1644
rect 4124 1636 4132 1644
rect 4460 1636 4468 1644
rect 4556 1636 4564 1644
rect 4812 1636 4820 1644
rect 4988 1636 4996 1644
rect 5468 1636 5476 1644
rect 1566 1606 1574 1614
rect 1580 1606 1588 1614
rect 1594 1606 1602 1614
rect 4638 1606 4646 1614
rect 4652 1606 4660 1614
rect 4666 1606 4674 1614
rect 876 1576 884 1584
rect 2316 1576 2324 1584
rect 2380 1576 2388 1584
rect 2460 1576 2468 1584
rect 2636 1576 2644 1584
rect 3196 1576 3204 1584
rect 3276 1576 3284 1584
rect 3452 1576 3460 1584
rect 5468 1576 5476 1584
rect 6236 1576 6244 1584
rect 1692 1556 1700 1564
rect 3020 1556 3028 1564
rect 892 1536 900 1544
rect 1100 1536 1108 1544
rect 1500 1536 1508 1544
rect 2300 1536 2308 1544
rect 2364 1536 2372 1544
rect 2444 1536 2452 1544
rect 2620 1536 2628 1544
rect 2780 1536 2788 1544
rect 2828 1536 2836 1544
rect 2860 1536 2868 1544
rect 3068 1536 3076 1544
rect 3868 1556 3876 1564
rect 4060 1556 4068 1564
rect 4108 1556 4116 1564
rect 4924 1556 4932 1564
rect 5692 1556 5700 1564
rect 3724 1536 3732 1544
rect 4092 1536 4100 1544
rect 4460 1536 4468 1544
rect 4860 1536 4868 1544
rect 4908 1536 4916 1544
rect 5100 1536 5108 1544
rect 5292 1536 5300 1544
rect 5708 1536 5716 1544
rect 12 1516 20 1524
rect 204 1516 212 1524
rect 428 1516 436 1524
rect 588 1516 596 1524
rect 812 1516 820 1524
rect 860 1516 868 1524
rect 1020 1516 1028 1524
rect 1036 1516 1044 1524
rect 1132 1516 1140 1524
rect 1196 1516 1204 1524
rect 92 1496 100 1504
rect 156 1496 164 1504
rect 268 1496 276 1504
rect 332 1496 340 1504
rect 348 1496 356 1504
rect 412 1496 420 1504
rect 476 1496 484 1504
rect 508 1496 516 1504
rect 556 1496 564 1504
rect 668 1496 676 1504
rect 796 1496 804 1504
rect 876 1496 884 1504
rect 988 1496 996 1504
rect 1084 1496 1092 1504
rect 1164 1496 1172 1504
rect 1244 1496 1252 1504
rect 1292 1496 1300 1504
rect 1772 1516 1780 1524
rect 1836 1516 1844 1524
rect 1932 1516 1940 1524
rect 2108 1516 2116 1524
rect 2332 1516 2340 1524
rect 2396 1516 2404 1524
rect 2412 1516 2420 1524
rect 2540 1516 2548 1524
rect 2588 1516 2596 1524
rect 2828 1516 2836 1524
rect 2892 1516 2900 1524
rect 2940 1516 2948 1524
rect 2956 1516 2964 1524
rect 3036 1516 3044 1524
rect 3100 1516 3108 1524
rect 3148 1516 3156 1524
rect 3260 1516 3268 1524
rect 3340 1516 3348 1524
rect 3420 1516 3428 1524
rect 3468 1516 3476 1524
rect 3548 1516 3556 1524
rect 3644 1516 3652 1524
rect 3788 1516 3796 1524
rect 3964 1516 3972 1524
rect 4028 1516 4036 1524
rect 4124 1516 4132 1524
rect 4172 1516 4180 1524
rect 4284 1516 4292 1524
rect 4332 1516 4340 1524
rect 4396 1516 4404 1524
rect 4492 1516 4500 1524
rect 4556 1516 4564 1524
rect 4572 1516 4580 1524
rect 4716 1516 4724 1524
rect 4828 1516 4836 1524
rect 4940 1516 4948 1524
rect 5068 1516 5076 1524
rect 5132 1516 5140 1524
rect 5324 1516 5332 1524
rect 5436 1516 5444 1524
rect 5708 1516 5716 1524
rect 5788 1516 5796 1524
rect 5836 1516 5844 1524
rect 5900 1516 5908 1524
rect 1340 1496 1348 1504
rect 1548 1496 1556 1504
rect 1724 1496 1732 1504
rect 1788 1496 1796 1504
rect 1852 1496 1860 1504
rect 44 1476 52 1484
rect 76 1476 84 1484
rect 124 1476 132 1484
rect 156 1476 164 1484
rect 252 1476 260 1484
rect 316 1476 324 1484
rect 364 1476 372 1484
rect 396 1476 404 1484
rect 460 1476 468 1484
rect 572 1476 580 1484
rect 620 1476 628 1484
rect 684 1476 692 1484
rect 700 1476 708 1484
rect 716 1480 724 1488
rect 2060 1496 2068 1504
rect 2188 1496 2196 1504
rect 2316 1496 2324 1504
rect 2380 1496 2388 1504
rect 2428 1496 2436 1504
rect 2636 1496 2644 1504
rect 2700 1496 2708 1504
rect 2764 1496 2772 1504
rect 2812 1496 2820 1504
rect 2876 1496 2884 1504
rect 2956 1496 2964 1504
rect 3084 1496 3092 1504
rect 3196 1496 3204 1504
rect 3308 1496 3316 1504
rect 3484 1496 3492 1504
rect 3612 1496 3620 1504
rect 3692 1496 3700 1504
rect 3756 1496 3764 1504
rect 3932 1496 3940 1504
rect 3948 1496 3956 1504
rect 3996 1496 4004 1504
rect 4108 1496 4116 1504
rect 4220 1496 4228 1504
rect 844 1476 852 1484
rect 956 1476 964 1484
rect 988 1476 996 1484
rect 1068 1476 1076 1484
rect 1084 1476 1092 1484
rect 1148 1476 1156 1484
rect 1260 1476 1268 1484
rect 1276 1476 1284 1484
rect 1356 1476 1364 1484
rect 204 1456 212 1464
rect 220 1456 228 1464
rect 284 1456 292 1464
rect 508 1456 516 1464
rect 764 1456 772 1464
rect 796 1456 804 1464
rect 924 1456 932 1464
rect 1372 1456 1380 1464
rect 1404 1476 1412 1484
rect 1436 1476 1444 1484
rect 1532 1476 1540 1484
rect 1596 1476 1604 1484
rect 1660 1476 1668 1484
rect 1708 1476 1716 1484
rect 1836 1476 1844 1484
rect 1900 1476 1908 1484
rect 1996 1476 2004 1484
rect 2012 1480 2020 1488
rect 2140 1476 2148 1484
rect 2492 1476 2500 1484
rect 2508 1476 2516 1484
rect 2556 1476 2564 1484
rect 2588 1476 2596 1484
rect 2716 1476 2724 1484
rect 2748 1476 2756 1484
rect 2908 1476 2916 1484
rect 3004 1476 3012 1484
rect 3212 1476 3220 1484
rect 3228 1476 3236 1484
rect 3340 1476 3348 1484
rect 3372 1476 3380 1484
rect 3388 1476 3396 1484
rect 3436 1476 3444 1484
rect 3516 1476 3524 1484
rect 3580 1476 3588 1484
rect 3596 1476 3604 1484
rect 3804 1476 3812 1484
rect 3900 1476 3908 1484
rect 3916 1476 3924 1484
rect 3980 1476 3988 1484
rect 4028 1476 4036 1484
rect 4140 1476 4148 1484
rect 4252 1496 4260 1504
rect 4364 1496 4372 1504
rect 4524 1496 4532 1504
rect 4540 1496 4548 1504
rect 4588 1496 4596 1504
rect 4812 1496 4820 1504
rect 4844 1496 4852 1504
rect 4876 1496 4884 1504
rect 4924 1496 4932 1504
rect 4956 1496 4964 1504
rect 5052 1496 5060 1504
rect 5100 1496 5108 1504
rect 5196 1496 5204 1504
rect 5308 1496 5316 1504
rect 5340 1496 5348 1504
rect 5468 1496 5476 1504
rect 5564 1496 5572 1504
rect 5692 1496 5700 1504
rect 5724 1496 5732 1504
rect 5852 1496 5860 1504
rect 5868 1496 5876 1504
rect 6140 1496 6148 1504
rect 4252 1476 4260 1484
rect 4284 1476 4292 1484
rect 4348 1476 4356 1484
rect 4444 1476 4452 1484
rect 4508 1476 4516 1484
rect 4636 1480 4644 1488
rect 4652 1476 4660 1484
rect 4748 1476 4756 1484
rect 4796 1476 4804 1484
rect 4972 1476 4980 1484
rect 5084 1476 5092 1484
rect 5180 1476 5188 1484
rect 5356 1476 5364 1484
rect 5404 1476 5412 1484
rect 5484 1476 5492 1484
rect 5580 1476 5588 1484
rect 5740 1476 5748 1484
rect 5788 1476 5796 1484
rect 5820 1476 5828 1484
rect 5884 1476 5892 1484
rect 5916 1476 5924 1484
rect 5932 1476 5940 1484
rect 5948 1476 5956 1484
rect 6044 1476 6052 1484
rect 6076 1476 6084 1484
rect 1404 1456 1412 1464
rect 1580 1456 1588 1464
rect 1644 1456 1652 1464
rect 1948 1456 1956 1464
rect 1980 1456 1988 1464
rect 2092 1456 2100 1464
rect 2156 1456 2164 1464
rect 2204 1456 2212 1464
rect 2236 1456 2244 1464
rect 2252 1456 2260 1464
rect 2476 1456 2484 1464
rect 2684 1456 2692 1464
rect 3660 1456 3668 1464
rect 4044 1456 4052 1464
rect 4412 1456 4420 1464
rect 4588 1456 4596 1464
rect 4668 1456 4676 1464
rect 4764 1456 4772 1464
rect 5004 1456 5012 1464
rect 5020 1456 5028 1464
rect 5052 1456 5060 1464
rect 5164 1456 5172 1464
rect 5388 1456 5396 1464
rect 5644 1456 5652 1464
rect 5772 1456 5780 1464
rect 12 1436 20 1444
rect 140 1436 148 1444
rect 236 1436 244 1444
rect 300 1436 308 1444
rect 364 1436 372 1444
rect 444 1436 452 1444
rect 492 1436 500 1444
rect 604 1436 612 1444
rect 636 1436 644 1444
rect 748 1436 756 1444
rect 780 1436 788 1444
rect 940 1436 948 1444
rect 1020 1436 1028 1444
rect 1052 1436 1060 1444
rect 1212 1436 1220 1444
rect 1324 1436 1332 1444
rect 1420 1436 1428 1444
rect 1964 1436 1972 1444
rect 2044 1436 2052 1444
rect 2076 1436 2084 1444
rect 2124 1436 2132 1444
rect 2268 1436 2276 1444
rect 2524 1436 2532 1444
rect 2636 1436 2644 1444
rect 2732 1436 2740 1444
rect 2860 1436 2868 1444
rect 2972 1436 2980 1444
rect 3244 1436 3252 1444
rect 3340 1436 3348 1444
rect 3420 1436 3428 1444
rect 3564 1436 3572 1444
rect 3644 1436 3652 1444
rect 3788 1436 3796 1444
rect 4172 1436 4180 1444
rect 4188 1436 4196 1444
rect 4284 1436 4292 1444
rect 4332 1436 4340 1444
rect 4396 1436 4404 1444
rect 4780 1436 4788 1444
rect 4988 1436 4996 1444
rect 5244 1436 5252 1444
rect 5308 1436 5316 1444
rect 5420 1436 5428 1444
rect 5580 1436 5588 1444
rect 5804 1436 5812 1444
rect 6012 1436 6020 1444
rect 3118 1406 3126 1414
rect 3132 1406 3140 1414
rect 3146 1406 3154 1414
rect 348 1376 356 1384
rect 876 1376 884 1384
rect 1068 1376 1076 1384
rect 1356 1376 1364 1384
rect 1916 1376 1924 1384
rect 2220 1376 2228 1384
rect 2428 1376 2436 1384
rect 2492 1376 2500 1384
rect 2652 1376 2660 1384
rect 2684 1376 2692 1384
rect 2764 1376 2772 1384
rect 3036 1376 3044 1384
rect 3260 1376 3268 1384
rect 3292 1376 3300 1384
rect 3804 1376 3812 1384
rect 3868 1376 3876 1384
rect 4204 1376 4212 1384
rect 5276 1376 5284 1384
rect 5436 1376 5444 1384
rect 5580 1376 5588 1384
rect 5756 1376 5764 1384
rect 5900 1376 5908 1384
rect 5932 1376 5940 1384
rect 12 1356 20 1364
rect 92 1356 100 1364
rect 620 1356 628 1364
rect 668 1356 676 1364
rect 748 1356 756 1364
rect 892 1356 900 1364
rect 924 1356 932 1364
rect 956 1356 964 1364
rect 1052 1356 1060 1364
rect 1372 1356 1380 1364
rect 1740 1356 1748 1364
rect 1772 1356 1780 1364
rect 1852 1356 1860 1364
rect 1932 1356 1940 1364
rect 1996 1356 2004 1364
rect 2108 1356 2116 1364
rect 2236 1356 2244 1364
rect 2396 1356 2404 1364
rect 2476 1356 2484 1364
rect 2668 1356 2676 1364
rect 2956 1356 2964 1364
rect 3084 1356 3092 1364
rect 3404 1356 3412 1364
rect 3452 1356 3460 1364
rect 3532 1356 3540 1364
rect 3948 1356 3956 1364
rect 3964 1356 3972 1364
rect 4076 1356 4084 1364
rect 4108 1356 4116 1364
rect 4140 1356 4148 1364
rect 4252 1356 4260 1364
rect 4268 1356 4276 1364
rect 4364 1356 4372 1364
rect 4812 1356 4820 1364
rect 4940 1356 4948 1364
rect 5196 1356 5204 1364
rect 5260 1356 5268 1364
rect 5420 1356 5428 1364
rect 5660 1356 5668 1364
rect 5756 1356 5764 1364
rect 5916 1356 5924 1364
rect 5996 1356 6004 1364
rect 300 1336 308 1344
rect 556 1336 564 1344
rect 636 1336 644 1344
rect 652 1336 660 1344
rect 716 1336 724 1344
rect 748 1336 756 1344
rect 812 1336 820 1344
rect 828 1336 836 1344
rect 956 1336 964 1344
rect 1036 1336 1044 1344
rect 1244 1336 1252 1344
rect 1276 1336 1284 1344
rect 1340 1336 1348 1344
rect 1452 1336 1460 1344
rect 1692 1336 1700 1344
rect 1772 1336 1780 1344
rect 1820 1336 1828 1344
rect 1884 1336 1892 1344
rect 1900 1336 1908 1344
rect 1948 1336 1956 1344
rect 2012 1336 2020 1344
rect 2092 1336 2100 1344
rect 2188 1336 2196 1344
rect 2204 1336 2212 1344
rect 2252 1336 2260 1344
rect 2508 1336 2516 1344
rect 2604 1336 2612 1344
rect 2700 1336 2708 1344
rect 2908 1336 2916 1344
rect 2972 1336 2980 1344
rect 3004 1336 3012 1344
rect 3068 1336 3076 1344
rect 3212 1336 3220 1344
rect 3276 1336 3284 1344
rect 3452 1336 3460 1344
rect 3612 1336 3620 1344
rect 3628 1336 3636 1344
rect 3692 1336 3700 1344
rect 3708 1336 3716 1344
rect 3772 1336 3780 1344
rect 3788 1336 3796 1344
rect 3916 1336 3924 1344
rect 3964 1336 3972 1344
rect 4012 1336 4020 1344
rect 4044 1336 4052 1344
rect 4156 1336 4164 1344
rect 4220 1336 4228 1344
rect 4284 1336 4292 1344
rect 4492 1336 4500 1344
rect 4540 1336 4548 1344
rect 4604 1336 4612 1344
rect 4636 1336 4644 1344
rect 4764 1336 4772 1344
rect 4828 1336 4836 1344
rect 4876 1336 4884 1344
rect 5004 1336 5012 1344
rect 5036 1336 5044 1344
rect 5132 1332 5140 1340
rect 5148 1336 5156 1344
rect 5212 1336 5220 1344
rect 5260 1336 5268 1344
rect 5292 1336 5300 1344
rect 5468 1336 5476 1344
rect 5628 1336 5636 1344
rect 5692 1336 5700 1344
rect 5756 1336 5764 1344
rect 5868 1336 5876 1344
rect 5948 1336 5956 1344
rect 6012 1336 6020 1344
rect 6076 1336 6084 1344
rect 44 1316 52 1324
rect 124 1316 132 1324
rect 204 1316 212 1324
rect 252 1316 260 1324
rect 316 1316 324 1324
rect 396 1316 404 1324
rect 460 1316 468 1324
rect 508 1316 516 1324
rect 524 1316 532 1324
rect 700 1316 708 1324
rect 780 1316 788 1324
rect 812 1316 820 1324
rect 844 1316 852 1324
rect 924 1316 932 1324
rect 972 1316 980 1324
rect 1084 1316 1092 1324
rect 1196 1316 1204 1324
rect 1228 1316 1236 1324
rect 1292 1316 1300 1324
rect 28 1296 36 1304
rect 108 1296 116 1304
rect 220 1296 228 1304
rect 236 1296 244 1304
rect 348 1296 356 1304
rect 412 1296 420 1304
rect 476 1296 484 1304
rect 492 1296 500 1304
rect 684 1296 692 1304
rect 764 1296 772 1304
rect 876 1296 884 1304
rect 1020 1296 1028 1304
rect 1212 1296 1220 1304
rect 1244 1296 1252 1304
rect 1468 1316 1476 1324
rect 1548 1316 1556 1324
rect 1660 1316 1668 1324
rect 1692 1316 1700 1324
rect 1788 1316 1796 1324
rect 1804 1316 1812 1324
rect 1884 1316 1892 1324
rect 1948 1316 1956 1324
rect 1980 1316 1988 1324
rect 2028 1316 2036 1324
rect 2060 1316 2068 1324
rect 2140 1316 2148 1324
rect 2188 1316 2196 1324
rect 2268 1316 2276 1324
rect 2300 1316 2308 1324
rect 2348 1316 2356 1324
rect 2444 1316 2452 1324
rect 2524 1316 2532 1324
rect 2556 1316 2564 1324
rect 2620 1316 2628 1324
rect 2716 1316 2724 1324
rect 2812 1316 2820 1324
rect 2860 1316 2868 1324
rect 2908 1316 2916 1324
rect 2940 1316 2948 1324
rect 2988 1316 2996 1324
rect 3020 1316 3028 1324
rect 1388 1296 1396 1304
rect 1500 1296 1508 1304
rect 1564 1296 1572 1304
rect 1676 1296 1684 1304
rect 1740 1296 1748 1304
rect 1836 1296 1844 1304
rect 2172 1296 2180 1304
rect 2316 1296 2324 1304
rect 2444 1296 2452 1304
rect 2540 1296 2548 1304
rect 2588 1296 2596 1304
rect 2764 1296 2772 1304
rect 2828 1296 2836 1304
rect 2844 1296 2852 1304
rect 3020 1296 3028 1304
rect 3180 1316 3188 1324
rect 3228 1316 3236 1324
rect 3356 1316 3364 1324
rect 3420 1316 3428 1324
rect 3484 1316 3492 1324
rect 3596 1316 3604 1324
rect 3644 1316 3652 1324
rect 3676 1316 3684 1324
rect 3724 1316 3732 1324
rect 3756 1316 3764 1324
rect 3868 1316 3876 1324
rect 3900 1316 3908 1324
rect 4028 1316 4036 1324
rect 4108 1316 4116 1324
rect 4156 1316 4164 1324
rect 4332 1316 4340 1324
rect 4412 1316 4420 1324
rect 4444 1316 4452 1324
rect 4540 1316 4548 1324
rect 4556 1316 4564 1324
rect 3196 1296 3204 1304
rect 3308 1296 3316 1304
rect 3468 1296 3476 1304
rect 3820 1296 3828 1304
rect 3884 1296 3892 1304
rect 4204 1296 4212 1304
rect 4252 1296 4260 1304
rect 108 1276 116 1284
rect 140 1276 148 1284
rect 268 1276 276 1284
rect 284 1276 292 1284
rect 380 1276 388 1284
rect 444 1276 452 1284
rect 1180 1276 1188 1284
rect 1324 1276 1332 1284
rect 1532 1276 1540 1284
rect 1644 1276 1652 1284
rect 2428 1276 2436 1284
rect 2572 1276 2580 1284
rect 2796 1276 2804 1284
rect 2876 1276 2884 1284
rect 3036 1276 3044 1284
rect 3340 1276 3348 1284
rect 3500 1276 3508 1284
rect 3644 1276 3652 1284
rect 3852 1276 3860 1284
rect 4316 1276 4324 1284
rect 4492 1296 4500 1304
rect 4524 1296 4532 1304
rect 4588 1296 4596 1304
rect 4716 1316 4724 1324
rect 4796 1316 4804 1324
rect 4892 1316 4900 1324
rect 5020 1316 5028 1324
rect 5052 1316 5060 1324
rect 5164 1316 5172 1324
rect 5292 1316 5300 1324
rect 5436 1316 5444 1324
rect 5580 1316 5588 1324
rect 5612 1316 5620 1324
rect 5772 1316 5780 1324
rect 5868 1316 5876 1324
rect 5964 1316 5972 1324
rect 6108 1318 6116 1326
rect 4764 1296 4772 1304
rect 4796 1296 4804 1304
rect 5084 1296 5092 1304
rect 5244 1296 5252 1304
rect 5340 1296 5348 1304
rect 5532 1296 5540 1304
rect 5596 1296 5604 1304
rect 5852 1296 5860 1304
rect 5900 1296 5908 1304
rect 6012 1296 6020 1304
rect 6044 1296 6052 1304
rect 4460 1276 4468 1284
rect 5500 1276 5508 1284
rect 5564 1276 5572 1284
rect 2028 1256 2036 1264
rect 2812 1256 2820 1264
rect 124 1236 132 1244
rect 204 1236 212 1244
rect 364 1236 372 1244
rect 460 1236 468 1244
rect 572 1236 580 1244
rect 940 1236 948 1244
rect 988 1236 996 1244
rect 1196 1236 1204 1244
rect 1420 1236 1428 1244
rect 1468 1236 1476 1244
rect 1516 1236 1524 1244
rect 1628 1236 1636 1244
rect 1756 1236 1764 1244
rect 2348 1236 2356 1244
rect 2860 1236 2868 1244
rect 3180 1236 3188 1244
rect 3356 1236 3364 1244
rect 3484 1236 3492 1244
rect 3548 1236 3556 1244
rect 3596 1236 3604 1244
rect 3756 1236 3764 1244
rect 4124 1236 4132 1244
rect 4348 1236 4356 1244
rect 4924 1236 4932 1244
rect 4972 1236 4980 1244
rect 5052 1236 5060 1244
rect 5100 1236 5108 1244
rect 5180 1236 5188 1244
rect 5324 1236 5332 1244
rect 6028 1236 6036 1244
rect 6236 1236 6244 1244
rect 1566 1206 1574 1214
rect 1580 1206 1588 1214
rect 1594 1206 1602 1214
rect 4638 1206 4646 1214
rect 4652 1206 4660 1214
rect 4666 1206 4674 1214
rect 492 1176 500 1184
rect 1452 1176 1460 1184
rect 1740 1176 1748 1184
rect 1820 1176 1828 1184
rect 1868 1176 1876 1184
rect 2076 1176 2084 1184
rect 2284 1176 2292 1184
rect 2332 1176 2340 1184
rect 2380 1176 2388 1184
rect 2476 1176 2484 1184
rect 2700 1176 2708 1184
rect 3164 1176 3172 1184
rect 3324 1176 3332 1184
rect 3708 1176 3716 1184
rect 3756 1176 3764 1184
rect 4012 1176 4020 1184
rect 4172 1176 4180 1184
rect 4204 1176 4212 1184
rect 4812 1176 4820 1184
rect 5244 1176 5252 1184
rect 1948 1156 1956 1164
rect 1436 1136 1444 1144
rect 1500 1136 1508 1144
rect 1804 1136 1812 1144
rect 1820 1136 1828 1144
rect 1932 1136 1940 1144
rect 1996 1136 2004 1144
rect 2140 1156 2148 1164
rect 2028 1136 2036 1144
rect 2060 1136 2068 1144
rect 2124 1136 2132 1144
rect 2188 1136 2196 1144
rect 3052 1156 3060 1164
rect 2220 1136 2228 1144
rect 2236 1136 2244 1144
rect 2316 1136 2324 1144
rect 2444 1136 2452 1144
rect 2572 1136 2580 1144
rect 2652 1136 2660 1144
rect 2924 1136 2932 1144
rect 3100 1136 3108 1144
rect 3196 1136 3204 1144
rect 3324 1136 3332 1144
rect 3340 1136 3348 1144
rect 3580 1136 3588 1144
rect 3692 1136 3700 1144
rect 4380 1136 4388 1144
rect 5372 1136 5380 1144
rect 5452 1136 5460 1144
rect 5596 1136 5604 1144
rect 188 1116 196 1124
rect 252 1116 260 1124
rect 348 1116 356 1124
rect 508 1116 516 1124
rect 620 1116 628 1124
rect 636 1116 644 1124
rect 700 1116 708 1124
rect 764 1116 772 1124
rect 812 1116 820 1124
rect 940 1116 948 1124
rect 1036 1116 1044 1124
rect 1116 1116 1124 1124
rect 1308 1116 1316 1124
rect 1468 1116 1476 1124
rect 1564 1116 1572 1124
rect 1708 1116 1716 1124
rect 1772 1116 1780 1124
rect 1820 1116 1828 1124
rect 1852 1116 1860 1124
rect 1964 1116 1972 1124
rect 2012 1116 2020 1124
rect 2092 1116 2100 1124
rect 2156 1116 2164 1124
rect 2220 1116 2228 1124
rect 2236 1116 2244 1124
rect 2348 1116 2356 1124
rect 2364 1116 2372 1124
rect 2428 1116 2436 1124
rect 2652 1116 2660 1124
rect 2684 1116 2692 1124
rect 2892 1116 2900 1124
rect 2956 1116 2964 1124
rect 3068 1116 3076 1124
rect 3228 1116 3236 1124
rect 3308 1116 3316 1124
rect 3372 1116 3380 1124
rect 3484 1116 3492 1124
rect 3516 1116 3524 1124
rect 3724 1116 3732 1124
rect 3948 1116 3956 1124
rect 4028 1116 4036 1124
rect 4252 1116 4260 1124
rect 4428 1116 4436 1124
rect 4716 1116 4724 1124
rect 4780 1116 4788 1124
rect 4828 1116 4836 1124
rect 4908 1116 4916 1124
rect 5228 1116 5236 1124
rect 5340 1116 5348 1124
rect 5484 1116 5492 1124
rect 5724 1116 5732 1124
rect 108 1096 116 1104
rect 156 1096 164 1104
rect 220 1096 228 1104
rect 268 1096 276 1104
rect 348 1096 356 1104
rect 396 1096 404 1104
rect 460 1096 468 1104
rect 524 1096 532 1104
rect 556 1096 564 1104
rect 668 1096 676 1104
rect 732 1096 740 1104
rect 860 1096 868 1104
rect 908 1096 916 1104
rect 972 1096 980 1104
rect 1068 1096 1076 1104
rect 1180 1096 1188 1104
rect 1260 1096 1268 1104
rect 1276 1096 1284 1104
rect 1308 1096 1316 1104
rect 1404 1096 1412 1104
rect 1452 1096 1460 1104
rect 1516 1096 1524 1104
rect 1596 1096 1604 1104
rect 1676 1096 1684 1104
rect 1724 1096 1732 1104
rect 1740 1096 1748 1104
rect 1820 1096 1828 1104
rect 1868 1096 1876 1104
rect 1948 1096 1956 1104
rect 2012 1096 2020 1104
rect 2076 1096 2084 1104
rect 2140 1096 2148 1104
rect 2204 1096 2212 1104
rect 2252 1096 2260 1104
rect 2332 1096 2340 1104
rect 2380 1096 2388 1104
rect 2444 1096 2452 1104
rect 2636 1096 2644 1104
rect 2668 1096 2676 1104
rect 2844 1096 2852 1104
rect 2876 1096 2884 1104
rect 2908 1096 2916 1104
rect 2988 1096 2996 1104
rect 3036 1096 3044 1104
rect 3084 1096 3092 1104
rect 3212 1096 3220 1104
rect 3244 1096 3252 1104
rect 3324 1096 3332 1104
rect 3436 1096 3444 1104
rect 3548 1096 3556 1104
rect 3596 1096 3604 1104
rect 3660 1096 3668 1104
rect 3708 1096 3716 1104
rect 3756 1096 3764 1104
rect 3836 1096 3844 1104
rect 3900 1096 3908 1104
rect 3996 1096 4004 1104
rect 4060 1096 4068 1104
rect 4108 1096 4116 1104
rect 4156 1096 4164 1104
rect 4252 1096 4260 1104
rect 4460 1096 4468 1104
rect 4556 1096 4564 1104
rect 4636 1096 4644 1104
rect 92 1076 100 1084
rect 108 1076 116 1084
rect 204 1076 212 1084
rect 268 1076 276 1084
rect 316 1076 324 1084
rect 380 1076 388 1084
rect 412 1076 420 1084
rect 444 1076 452 1084
rect 572 1076 580 1084
rect 588 1076 596 1084
rect 684 1076 692 1084
rect 748 1076 756 1084
rect 796 1076 804 1084
rect 844 1076 852 1084
rect 860 1076 868 1084
rect 924 1076 932 1084
rect 972 1076 980 1084
rect 988 1076 996 1084
rect 1020 1076 1028 1084
rect 1052 1076 1060 1084
rect 1164 1076 1172 1084
rect 1260 1076 1268 1084
rect 1292 1076 1300 1084
rect 1372 1076 1380 1084
rect 1404 1076 1412 1084
rect 1612 1076 1620 1084
rect 1660 1076 1668 1084
rect 1724 1076 1732 1084
rect 2508 1076 2516 1084
rect 2620 1076 2628 1084
rect 2764 1076 2772 1084
rect 2796 1076 2804 1084
rect 2908 1076 2916 1084
rect 2972 1076 2980 1084
rect 3212 1076 3220 1084
rect 3260 1076 3268 1084
rect 3404 1076 3412 1084
rect 3420 1076 3428 1084
rect 3452 1076 3460 1084
rect 3484 1076 3492 1084
rect 3532 1076 3540 1084
rect 3612 1076 3620 1084
rect 3644 1076 3652 1084
rect 3740 1076 3748 1084
rect 3820 1076 3828 1084
rect 3980 1076 3988 1084
rect 4076 1076 4084 1084
rect 4092 1076 4100 1084
rect 4220 1076 4228 1084
rect 4284 1076 4292 1084
rect 4412 1076 4420 1084
rect 4476 1076 4484 1084
rect 4492 1076 4500 1084
rect 4588 1076 4596 1084
rect 4956 1096 4964 1104
rect 5196 1096 5204 1104
rect 5228 1096 5236 1104
rect 5276 1096 5284 1104
rect 5356 1096 5364 1104
rect 5580 1096 5588 1104
rect 5660 1096 5668 1104
rect 5708 1096 5716 1104
rect 5740 1096 5748 1104
rect 5788 1096 5796 1104
rect 108 1056 116 1064
rect 1244 1056 1252 1064
rect 1340 1056 1348 1064
rect 1356 1056 1364 1064
rect 1644 1056 1652 1064
rect 2540 1056 2548 1064
rect 2556 1056 2564 1064
rect 2588 1056 2596 1064
rect 2780 1056 2788 1064
rect 3036 1056 3044 1064
rect 3292 1056 3300 1064
rect 3372 1056 3380 1064
rect 3644 1056 3652 1064
rect 3820 1056 3828 1064
rect 3900 1056 3908 1064
rect 3932 1056 3940 1064
rect 3996 1056 4004 1064
rect 4156 1056 4164 1064
rect 4188 1056 4196 1064
rect 4268 1056 4276 1064
rect 4300 1056 4308 1064
rect 4748 1076 4756 1084
rect 4860 1076 4868 1084
rect 4892 1076 4900 1084
rect 4940 1076 4948 1084
rect 5004 1076 5012 1084
rect 5100 1076 5108 1084
rect 5292 1076 5300 1084
rect 5404 1076 5412 1084
rect 5436 1076 5444 1084
rect 5916 1094 5924 1102
rect 6108 1094 6116 1102
rect 5852 1076 5860 1084
rect 5980 1076 5988 1084
rect 6076 1076 6084 1084
rect 4732 1056 4740 1064
rect 4844 1056 4852 1064
rect 4988 1056 4996 1064
rect 5132 1056 5140 1064
rect 5148 1056 5156 1064
rect 5260 1056 5268 1064
rect 5324 1056 5332 1064
rect 5404 1056 5412 1064
rect 5516 1056 5524 1064
rect 5532 1056 5540 1064
rect 5628 1056 5636 1064
rect 5676 1056 5684 1064
rect 5708 1056 5716 1064
rect 5916 1056 5924 1064
rect 92 1036 100 1044
rect 188 1036 196 1044
rect 284 1036 292 1044
rect 348 1036 356 1044
rect 428 1036 436 1044
rect 604 1036 612 1044
rect 636 1036 644 1044
rect 700 1036 708 1044
rect 780 1036 788 1044
rect 812 1036 820 1044
rect 908 1036 916 1044
rect 940 1036 948 1044
rect 1100 1036 1108 1044
rect 1116 1036 1124 1044
rect 1212 1036 1220 1044
rect 1516 1036 1524 1044
rect 2524 1036 2532 1044
rect 2604 1036 2612 1044
rect 3132 1036 3140 1044
rect 3164 1036 3172 1044
rect 3500 1036 3508 1044
rect 3868 1036 3876 1044
rect 3916 1036 3924 1044
rect 4028 1036 4036 1044
rect 4428 1036 4436 1044
rect 4908 1036 4916 1044
rect 4972 1036 4980 1044
rect 5068 1036 5076 1044
rect 5116 1036 5124 1044
rect 5244 1036 5252 1044
rect 5308 1036 5316 1044
rect 5500 1036 5508 1044
rect 5548 1036 5556 1044
rect 5580 1036 5588 1044
rect 5644 1036 5652 1044
rect 6044 1036 6052 1044
rect 6236 1036 6244 1044
rect 3118 1006 3126 1014
rect 3132 1006 3140 1014
rect 3146 1006 3154 1014
rect 156 976 164 984
rect 1884 976 1892 984
rect 1948 976 1956 984
rect 2140 976 2148 984
rect 2332 976 2340 984
rect 2908 976 2916 984
rect 2988 976 2996 984
rect 3100 976 3108 984
rect 3276 976 3284 984
rect 4060 976 4068 984
rect 4300 976 4308 984
rect 4364 976 4372 984
rect 4540 976 4548 984
rect 4988 976 4996 984
rect 5036 976 5044 984
rect 5276 976 5284 984
rect 5484 976 5492 984
rect 5548 976 5556 984
rect 6172 976 6180 984
rect 140 956 148 964
rect 380 956 388 964
rect 668 956 676 964
rect 748 956 756 964
rect 844 956 852 964
rect 940 956 948 964
rect 1068 956 1076 964
rect 1164 956 1172 964
rect 1324 956 1332 964
rect 1500 956 1508 964
rect 1772 956 1780 964
rect 2028 956 2036 964
rect 2076 956 2084 964
rect 2508 956 2516 964
rect 2620 956 2628 964
rect 2700 956 2708 964
rect 2860 956 2868 964
rect 3036 956 3044 964
rect 3388 956 3396 964
rect 3548 956 3556 964
rect 188 936 196 944
rect 332 936 340 944
rect 700 936 708 944
rect 732 936 740 944
rect 764 936 772 944
rect 1020 936 1028 944
rect 1196 936 1204 944
rect 1308 936 1316 944
rect 1564 936 1572 944
rect 1628 936 1636 944
rect 1724 936 1732 944
rect 1740 936 1748 944
rect 1836 936 1844 944
rect 1996 936 2004 944
rect 2044 936 2052 944
rect 2092 936 2100 944
rect 2284 936 2292 944
rect 2428 936 2436 944
rect 2460 936 2468 944
rect 2636 936 2644 944
rect 2716 936 2724 944
rect 2860 936 2868 944
rect 3020 936 3028 944
rect 3116 936 3124 944
rect 3228 936 3236 944
rect 3292 936 3300 944
rect 3372 936 3380 944
rect 3436 936 3444 944
rect 3452 936 3460 944
rect 3516 936 3524 944
rect 3564 936 3572 944
rect 3692 956 3700 964
rect 3708 956 3716 964
rect 3820 956 3828 964
rect 3852 956 3860 964
rect 4124 956 4132 964
rect 4220 956 4228 964
rect 4396 956 4404 964
rect 4460 956 4468 964
rect 4524 956 4532 964
rect 4588 956 4596 964
rect 4620 956 4628 964
rect 4700 956 4708 964
rect 4796 956 4804 964
rect 5052 956 5060 964
rect 3676 936 3684 944
rect 3868 936 3876 944
rect 3916 936 3924 944
rect 4044 936 4052 944
rect 4236 936 4244 944
rect 4332 936 4340 944
rect 4380 936 4388 944
rect 4428 936 4436 944
rect 4476 936 4484 944
rect 4524 936 4532 944
rect 4556 936 4564 944
rect 4588 936 4596 944
rect 4748 936 4756 944
rect 4844 936 4852 944
rect 4876 936 4884 944
rect 4892 936 4900 944
rect 4924 936 4932 944
rect 5020 936 5028 944
rect 5132 936 5140 944
rect 5196 936 5204 944
rect 5244 936 5252 944
rect 5340 936 5348 944
rect 5404 936 5412 944
rect 5580 956 5588 964
rect 5708 956 5716 964
rect 5516 936 5524 944
rect 5676 936 5684 944
rect 5788 956 5796 964
rect 6156 956 6164 964
rect 5996 936 6004 944
rect 6092 936 6100 944
rect 6236 936 6244 944
rect 44 916 52 924
rect 108 916 116 924
rect 188 916 196 924
rect 236 916 244 924
rect 300 916 308 924
rect 332 916 340 924
rect 428 916 436 924
rect 492 916 500 924
rect 540 916 548 924
rect 620 916 628 924
rect 716 916 724 924
rect 812 916 820 924
rect 892 916 900 924
rect 972 916 980 924
rect 1132 916 1140 924
rect 1228 916 1236 924
rect 60 896 68 904
rect 124 896 132 904
rect 252 896 260 904
rect 268 896 276 904
rect 444 896 452 904
rect 524 896 532 904
rect 620 896 628 904
rect 684 896 692 904
rect 908 896 916 904
rect 940 896 948 904
rect 1068 896 1076 904
rect 1148 896 1156 904
rect 1260 896 1268 904
rect 1388 916 1396 924
rect 1436 916 1444 924
rect 1612 916 1620 924
rect 1404 896 1412 904
rect 1420 896 1428 904
rect 1548 896 1556 904
rect 1660 896 1668 904
rect 1724 916 1732 924
rect 1804 916 1812 924
rect 1884 916 1892 924
rect 1948 916 1956 924
rect 1980 916 1988 924
rect 2028 916 2036 924
rect 2108 916 2116 924
rect 2188 916 2196 924
rect 2300 916 2308 924
rect 2380 916 2388 924
rect 2412 916 2420 924
rect 2476 916 2484 924
rect 2508 916 2516 924
rect 2540 916 2548 924
rect 2588 916 2596 924
rect 2652 916 2660 924
rect 2796 916 2804 924
rect 2828 916 2836 924
rect 3212 916 3220 924
rect 3276 916 3284 924
rect 3404 916 3412 924
rect 3468 916 3476 924
rect 3580 916 3588 924
rect 3612 916 3620 924
rect 3660 916 3668 924
rect 3788 916 3796 924
rect 3932 916 3940 924
rect 3996 916 4004 924
rect 4028 916 4036 924
rect 4092 916 4100 924
rect 4156 916 4164 924
rect 4172 916 4180 924
rect 4460 916 4468 924
rect 4572 916 4580 924
rect 4684 916 4692 924
rect 4732 916 4740 924
rect 4908 916 4916 924
rect 4956 916 4964 924
rect 5004 916 5012 924
rect 5100 916 5108 924
rect 5148 916 5156 924
rect 5164 916 5172 924
rect 5388 916 5396 924
rect 5452 916 5460 924
rect 5468 916 5476 924
rect 5628 916 5636 924
rect 5660 916 5668 924
rect 5740 916 5748 924
rect 5852 918 5860 926
rect 5916 916 5924 924
rect 6092 916 6100 924
rect 6188 916 6196 924
rect 6204 916 6212 924
rect 1788 896 1796 904
rect 1884 896 1892 904
rect 1964 896 1972 904
rect 2092 896 2100 904
rect 2204 896 2212 904
rect 2220 896 2228 904
rect 2332 896 2340 904
rect 2396 896 2404 904
rect 2540 896 2548 904
rect 2684 896 2692 904
rect 28 876 36 884
rect 92 876 100 884
rect 220 876 228 884
rect 284 876 292 884
rect 412 876 420 884
rect 476 876 484 884
rect 556 876 564 884
rect 604 876 612 884
rect 988 876 996 884
rect 1020 876 1028 884
rect 1084 876 1092 884
rect 1116 876 1124 884
rect 1340 876 1348 884
rect 1372 876 1380 884
rect 1436 876 1444 884
rect 1452 876 1460 884
rect 1820 876 1828 884
rect 1868 876 1876 884
rect 1948 876 1956 884
rect 2172 876 2180 884
rect 2396 876 2404 884
rect 2556 876 2564 884
rect 2588 876 2596 884
rect 2652 876 2660 884
rect 2780 876 2788 884
rect 2908 896 2916 904
rect 3292 896 3300 904
rect 3404 896 3412 904
rect 3500 896 3508 904
rect 3804 896 3812 904
rect 3948 896 3956 904
rect 4012 896 4020 904
rect 4348 896 4356 904
rect 4508 896 4516 904
rect 4796 896 4804 904
rect 4844 896 4852 904
rect 4860 896 4868 904
rect 4924 896 4932 904
rect 5116 896 5124 904
rect 5180 896 5188 904
rect 5212 896 5220 904
rect 5228 896 5236 904
rect 5356 896 5364 904
rect 5548 896 5556 904
rect 5644 896 5652 904
rect 3740 876 3748 884
rect 3772 876 3780 884
rect 3916 876 3924 884
rect 3980 876 3988 884
rect 4732 876 4740 884
rect 5084 876 5092 884
rect 5388 876 5396 884
rect 5612 876 5620 884
rect 5980 876 5988 884
rect 6140 876 6148 884
rect 1388 856 1396 864
rect 1484 856 1492 864
rect 1692 856 1700 864
rect 2188 856 2196 864
rect 2748 856 2756 864
rect 5100 856 5108 864
rect 5628 856 5636 864
rect 44 836 52 844
rect 108 836 116 844
rect 236 836 244 844
rect 284 836 292 844
rect 380 836 388 844
rect 428 836 436 844
rect 492 836 500 844
rect 540 836 548 844
rect 620 836 628 844
rect 796 836 804 844
rect 828 836 836 844
rect 892 836 900 844
rect 924 836 932 844
rect 972 836 980 844
rect 1132 836 1140 844
rect 1164 836 1172 844
rect 1292 836 1300 844
rect 1436 836 1444 844
rect 1772 836 1780 844
rect 2252 836 2260 844
rect 2380 836 2388 844
rect 2428 836 2436 844
rect 2492 836 2500 844
rect 2572 836 2580 844
rect 2764 836 2772 844
rect 2844 836 2852 844
rect 3180 836 3188 844
rect 3788 836 3796 844
rect 3836 836 3844 844
rect 3996 836 4004 844
rect 4604 836 4612 844
rect 5452 836 5460 844
rect 5564 836 5572 844
rect 6028 836 6036 844
rect 1566 806 1574 814
rect 1580 806 1588 814
rect 1594 806 1602 814
rect 4638 806 4646 814
rect 4652 806 4660 814
rect 4666 806 4674 814
rect 652 776 660 784
rect 1516 776 1524 784
rect 1548 776 1556 784
rect 1660 776 1668 784
rect 1836 776 1844 784
rect 1900 776 1908 784
rect 1948 776 1956 784
rect 1980 776 1988 784
rect 2028 776 2036 784
rect 2108 776 2116 784
rect 2188 776 2196 784
rect 2860 776 2868 784
rect 2924 776 2932 784
rect 3804 776 3812 784
rect 4460 776 4468 784
rect 4844 776 4852 784
rect 5052 776 5060 784
rect 6204 776 6212 784
rect 316 756 324 764
rect 2796 756 2804 764
rect 3724 756 3732 764
rect 5340 756 5348 764
rect 364 736 372 744
rect 412 736 420 744
rect 1564 736 1572 744
rect 1820 736 1828 744
rect 1884 736 1892 744
rect 1964 736 1972 744
rect 2012 736 2020 744
rect 2092 736 2100 744
rect 2140 736 2148 744
rect 2444 736 2452 744
rect 2812 736 2820 744
rect 2908 736 2916 744
rect 3308 736 3316 744
rect 3676 736 3684 744
rect 3708 736 3716 744
rect 4012 736 4020 744
rect 4700 736 4708 744
rect 4748 736 4756 744
rect 4780 736 4788 744
rect 4972 736 4980 744
rect 5324 736 5332 744
rect 5564 736 5572 744
rect 5772 736 5780 744
rect 6124 736 6132 744
rect 140 716 148 724
rect 252 716 260 724
rect 332 716 340 724
rect 380 716 388 724
rect 444 716 452 724
rect 460 716 468 724
rect 524 716 532 724
rect 588 716 596 724
rect 684 716 692 724
rect 780 716 788 724
rect 892 716 900 724
rect 940 716 948 724
rect 972 716 980 724
rect 1068 716 1076 724
rect 1100 716 1108 724
rect 1116 716 1124 724
rect 1228 716 1236 724
rect 1324 716 1332 724
rect 1532 716 1540 724
rect 1852 716 1860 724
rect 1916 716 1924 724
rect 2060 716 2068 724
rect 2236 716 2244 724
rect 2316 716 2324 724
rect 2364 716 2372 724
rect 2412 716 2420 724
rect 2476 716 2484 724
rect 2764 716 2772 724
rect 2780 716 2788 724
rect 2844 716 2852 724
rect 2940 716 2948 724
rect 3276 716 3284 724
rect 3404 716 3412 724
rect 3436 716 3444 724
rect 3500 716 3508 724
rect 3644 716 3652 724
rect 3740 716 3748 724
rect 3900 716 3908 724
rect 3916 716 3924 724
rect 4284 716 4292 724
rect 4364 716 4372 724
rect 4444 716 4452 724
rect 4476 716 4484 724
rect 4668 716 4676 724
rect 4812 716 4820 724
rect 4908 716 4916 724
rect 5004 716 5012 724
rect 5020 716 5028 724
rect 5116 716 5124 724
rect 5292 716 5300 724
rect 5356 716 5364 724
rect 5436 716 5444 724
rect 5532 716 5540 724
rect 6236 716 6244 724
rect 76 696 84 704
rect 172 696 180 704
rect 268 696 276 704
rect 348 696 356 704
rect 396 696 404 704
rect 508 696 516 704
rect 572 696 580 704
rect 652 696 660 704
rect 764 696 772 704
rect 844 696 852 704
rect 892 696 900 704
rect 92 676 100 684
rect 204 676 212 684
rect 236 676 244 684
rect 284 676 292 684
rect 396 676 404 684
rect 492 676 500 684
rect 524 676 532 684
rect 588 676 596 684
rect 620 676 628 684
rect 636 676 644 684
rect 716 676 724 684
rect 780 676 788 684
rect 812 676 820 684
rect 828 676 836 684
rect 924 676 932 684
rect 988 696 996 704
rect 1068 696 1076 704
rect 1148 696 1156 704
rect 1180 696 1188 704
rect 1260 696 1268 704
rect 1372 696 1380 704
rect 1468 696 1476 704
rect 1548 696 1556 704
rect 1836 696 1844 704
rect 1900 696 1908 704
rect 1948 696 1956 704
rect 2028 696 2036 704
rect 2076 696 2084 704
rect 2156 696 2164 704
rect 2172 696 2180 704
rect 2220 696 2228 704
rect 2284 696 2292 704
rect 2332 696 2340 704
rect 2460 696 2468 704
rect 2492 696 2500 704
rect 2652 696 2660 704
rect 2796 696 2804 704
rect 2924 696 2932 704
rect 2972 696 2980 704
rect 3020 696 3028 704
rect 3052 696 3060 704
rect 3068 696 3076 704
rect 3164 696 3172 704
rect 3212 696 3220 704
rect 3292 696 3300 704
rect 3340 696 3348 704
rect 3468 696 3476 704
rect 3548 696 3556 704
rect 3564 696 3572 704
rect 3660 696 3668 704
rect 3724 696 3732 704
rect 3916 696 3924 704
rect 3980 696 3988 704
rect 4156 696 4164 704
rect 4252 696 4260 704
rect 4364 696 4372 704
rect 4476 696 4484 704
rect 4540 696 4548 704
rect 4556 696 4564 704
rect 4684 696 4692 704
rect 4732 696 4740 704
rect 4796 696 4804 704
rect 4828 696 4836 704
rect 4876 696 4884 704
rect 5052 696 5060 704
rect 5196 696 5204 704
rect 5292 696 5300 704
rect 5340 696 5348 704
rect 5372 696 5380 704
rect 5516 696 5524 704
rect 5548 696 5556 704
rect 5660 696 5668 704
rect 5708 696 5716 704
rect 5820 696 5828 704
rect 5884 696 5892 704
rect 6028 696 6036 704
rect 6140 696 6148 704
rect 6204 696 6212 704
rect 988 676 996 684
rect 1036 676 1044 684
rect 1164 676 1172 684
rect 1276 676 1284 684
rect 1292 676 1300 684
rect 1388 676 1396 684
rect 1452 676 1460 684
rect 1708 676 1716 684
rect 76 656 84 664
rect 316 656 324 664
rect 588 656 596 664
rect 780 656 788 664
rect 1212 656 1220 664
rect 1340 656 1348 664
rect 1452 656 1460 664
rect 1516 656 1524 664
rect 1692 656 1700 664
rect 2124 656 2132 664
rect 2204 656 2212 664
rect 2268 676 2276 684
rect 2332 676 2340 684
rect 2364 676 2372 684
rect 2380 676 2388 684
rect 2508 676 2516 684
rect 2668 676 2676 684
rect 2876 676 2884 684
rect 2956 676 2964 684
rect 3068 676 3076 684
rect 3196 676 3204 684
rect 3260 676 3268 684
rect 3356 676 3364 684
rect 3388 676 3396 684
rect 3452 676 3460 684
rect 3484 676 3492 684
rect 3596 676 3604 684
rect 3772 676 3780 684
rect 3852 676 3860 684
rect 3948 676 3956 684
rect 3964 676 3972 684
rect 4028 676 4036 684
rect 4124 676 4132 684
rect 4140 676 4148 684
rect 4268 676 4276 684
rect 4332 676 4340 684
rect 4396 676 4404 684
rect 4444 676 4452 684
rect 4492 676 4500 684
rect 4572 676 4580 684
rect 4796 676 4804 684
rect 4956 676 4964 684
rect 5068 676 5076 684
rect 5084 676 5092 684
rect 5212 676 5220 684
rect 5260 676 5268 684
rect 5452 676 5460 684
rect 5468 676 5476 684
rect 5500 676 5508 684
rect 5788 676 5796 684
rect 5884 676 5892 684
rect 6172 676 6180 684
rect 6188 676 6196 684
rect 2540 656 2548 664
rect 2556 656 2564 664
rect 2604 656 2612 664
rect 2668 656 2676 664
rect 2700 656 2708 664
rect 2828 656 2836 664
rect 3020 656 3028 664
rect 3196 656 3204 664
rect 3260 656 3268 664
rect 3388 656 3396 664
rect 3516 656 3524 664
rect 3580 656 3588 664
rect 3660 656 3668 664
rect 3804 656 3812 664
rect 3820 656 3828 664
rect 4204 656 4212 664
rect 4300 656 4308 664
rect 4380 656 4388 664
rect 4540 656 4548 664
rect 4588 656 4596 664
rect 4604 656 4612 664
rect 4732 656 4740 664
rect 4828 656 4836 664
rect 4924 656 4932 664
rect 5228 656 5236 664
rect 5372 656 5380 664
rect 5996 656 6004 664
rect 92 636 100 644
rect 124 636 132 644
rect 252 636 260 644
rect 444 636 452 644
rect 460 636 468 644
rect 732 636 740 644
rect 908 636 916 644
rect 956 636 964 644
rect 1116 636 1124 644
rect 1228 636 1236 644
rect 1324 636 1332 644
rect 1404 636 1412 644
rect 1772 636 1780 644
rect 2140 636 2148 644
rect 2396 636 2404 644
rect 2444 636 2452 644
rect 2524 636 2532 644
rect 2668 636 2676 644
rect 2764 636 2772 644
rect 3292 636 3300 644
rect 3532 636 3540 644
rect 3916 636 3924 644
rect 4092 636 4100 644
rect 4188 636 4196 644
rect 4316 636 4324 644
rect 4908 636 4916 644
rect 5100 636 5108 644
rect 5180 636 5188 644
rect 5500 636 5508 644
rect 5580 636 5588 644
rect 5932 636 5940 644
rect 3118 606 3126 614
rect 3132 606 3140 614
rect 3146 606 3154 614
rect 60 576 68 584
rect 332 576 340 584
rect 668 576 676 584
rect 828 576 836 584
rect 1212 576 1220 584
rect 1356 576 1364 584
rect 1420 576 1428 584
rect 1596 576 1604 584
rect 1676 576 1684 584
rect 1740 576 1748 584
rect 1804 576 1812 584
rect 1868 576 1876 584
rect 1932 576 1940 584
rect 2044 576 2052 584
rect 2108 576 2116 584
rect 2156 576 2164 584
rect 2252 576 2260 584
rect 2348 576 2356 584
rect 2412 576 2420 584
rect 2476 576 2484 584
rect 2684 576 2692 584
rect 2748 576 2756 584
rect 3436 576 3444 584
rect 3580 576 3588 584
rect 3708 576 3716 584
rect 4284 576 4292 584
rect 4396 576 4404 584
rect 4780 576 4788 584
rect 4876 576 4884 584
rect 4972 576 4980 584
rect 6220 576 6228 584
rect 108 556 116 564
rect 140 556 148 564
rect 572 556 580 564
rect 652 556 660 564
rect 1164 556 1172 564
rect 1452 556 1460 564
rect 1628 556 1636 564
rect 1820 556 1828 564
rect 1884 556 1892 564
rect 2060 556 2068 564
rect 2124 556 2132 564
rect 2140 556 2148 564
rect 2604 556 2612 564
rect 2844 556 2852 564
rect 2876 556 2884 564
rect 3244 556 3252 564
rect 3276 556 3284 564
rect 3708 556 3716 564
rect 92 536 100 544
rect 188 536 196 544
rect 380 536 388 544
rect 540 536 548 544
rect 684 536 692 544
rect 732 536 740 544
rect 764 536 772 544
rect 892 536 900 544
rect 220 516 228 524
rect 300 516 308 524
rect 364 516 372 524
rect 492 516 500 524
rect 524 516 532 524
rect 572 516 580 524
rect 620 516 628 524
rect 700 516 708 524
rect 748 516 756 524
rect 860 516 868 524
rect 876 516 884 524
rect 1228 536 1236 544
rect 1308 536 1316 544
rect 1484 536 1492 544
rect 1788 536 1796 544
rect 1852 536 1860 544
rect 1996 536 2004 544
rect 2028 536 2036 544
rect 2092 536 2100 544
rect 2172 536 2180 544
rect 2236 536 2244 544
rect 2284 536 2292 544
rect 2380 536 2388 544
rect 2396 536 2404 544
rect 2444 536 2452 544
rect 2572 536 2580 544
rect 2604 536 2612 544
rect 2620 536 2628 544
rect 2716 536 2724 544
rect 2732 536 2740 544
rect 2780 536 2788 544
rect 2860 536 2868 544
rect 3020 536 3028 544
rect 3036 536 3044 544
rect 3116 536 3124 544
rect 3212 536 3220 544
rect 3244 536 3252 544
rect 3260 536 3268 544
rect 3308 536 3316 544
rect 3404 536 3412 544
rect 3420 536 3428 544
rect 3500 536 3508 544
rect 3516 536 3524 544
rect 3612 536 3620 544
rect 3724 536 3732 544
rect 3932 556 3940 564
rect 4412 556 4420 564
rect 4620 556 4628 564
rect 4716 556 4724 564
rect 4844 556 4852 564
rect 4860 556 4868 564
rect 4956 556 4964 564
rect 3804 536 3812 544
rect 3820 536 3828 544
rect 3884 536 3892 544
rect 3900 536 3908 544
rect 3932 536 3940 544
rect 4076 536 4084 544
rect 4156 536 4164 544
rect 4236 536 4244 544
rect 4380 536 4388 544
rect 4540 536 4548 544
rect 4588 536 4596 544
rect 4636 536 4644 544
rect 4812 536 4820 544
rect 4844 536 4852 544
rect 4972 536 4980 544
rect 5068 556 5076 564
rect 5084 556 5092 564
rect 5212 556 5220 564
rect 5308 556 5316 564
rect 5404 556 5412 564
rect 5676 556 5684 564
rect 5692 556 5700 564
rect 5852 556 5860 564
rect 5884 556 5892 564
rect 5916 556 5924 564
rect 5116 536 5124 544
rect 5244 536 5252 544
rect 5340 536 5348 544
rect 5468 536 5476 544
rect 5644 536 5652 544
rect 5756 536 5764 544
rect 5788 536 5796 544
rect 5980 536 5988 544
rect 5996 536 6004 544
rect 6252 536 6260 544
rect 924 516 932 524
rect 1004 516 1012 524
rect 1068 516 1076 524
rect 1116 516 1124 524
rect 1244 516 1252 524
rect 1276 516 1284 524
rect 1356 516 1364 524
rect 1404 516 1412 524
rect 1468 516 1476 524
rect 1500 516 1508 524
rect 1612 516 1620 524
rect 1676 516 1684 524
rect 1740 516 1748 524
rect 1772 516 1780 524
rect 1836 516 1844 524
rect 1916 516 1924 524
rect 2012 516 2020 524
rect 2076 516 2084 524
rect 2188 516 2196 524
rect 2220 516 2228 524
rect 2524 516 2532 524
rect 2556 516 2564 524
rect 2796 516 2804 524
rect 204 496 212 504
rect 316 496 324 504
rect 332 496 340 504
rect 444 496 452 504
rect 508 496 516 504
rect 636 496 644 504
rect 716 496 724 504
rect 828 496 836 504
rect 844 496 852 504
rect 956 496 964 504
rect 1020 496 1028 504
rect 1084 496 1092 504
rect 1164 496 1172 504
rect 1260 496 1268 504
rect 1372 496 1380 504
rect 140 476 148 484
rect 236 476 244 484
rect 284 476 292 484
rect 412 476 420 484
rect 476 476 484 484
rect 604 476 612 484
rect 988 476 996 484
rect 1052 476 1060 484
rect 1132 476 1140 484
rect 1292 476 1300 484
rect 1340 476 1348 484
rect 1356 476 1364 484
rect 1548 496 1556 504
rect 1692 496 1700 504
rect 1756 496 1764 504
rect 1900 496 1908 504
rect 1964 496 1972 504
rect 2220 496 2228 504
rect 2268 496 2276 504
rect 2428 496 2436 504
rect 2540 496 2548 504
rect 2764 496 2772 504
rect 2876 516 2884 524
rect 2892 516 2900 524
rect 2940 516 2948 524
rect 3004 516 3012 524
rect 3164 516 3172 524
rect 3196 516 3204 524
rect 3068 496 3076 504
rect 3180 496 3188 504
rect 3292 496 3300 504
rect 3372 496 3380 504
rect 3692 516 3700 524
rect 3468 496 3476 504
rect 3836 516 3844 524
rect 3868 516 3876 524
rect 3964 516 3972 524
rect 4028 516 4036 524
rect 4124 516 4132 524
rect 4188 516 4196 524
rect 4252 516 4260 524
rect 4316 516 4324 524
rect 4364 516 4372 524
rect 4444 516 4452 524
rect 4508 516 4516 524
rect 4748 516 4756 524
rect 4796 516 4804 524
rect 4956 516 4964 524
rect 5100 516 5108 524
rect 5132 516 5140 524
rect 5164 516 5172 524
rect 5356 516 5364 524
rect 5388 516 5396 524
rect 5420 516 5428 524
rect 5484 516 5492 524
rect 5516 516 5524 524
rect 5580 516 5588 524
rect 5628 516 5636 524
rect 5692 516 5700 524
rect 5740 516 5748 524
rect 5804 516 5812 524
rect 5820 516 5828 524
rect 6028 516 6036 524
rect 6124 516 6132 524
rect 6172 516 6180 524
rect 3868 496 3876 504
rect 3948 496 3956 504
rect 4012 496 4020 504
rect 4108 496 4116 504
rect 4220 496 4228 504
rect 4300 496 4308 504
rect 4348 496 4356 504
rect 4428 496 4436 504
rect 4492 496 4500 504
rect 4556 496 4564 504
rect 4716 496 4724 504
rect 5068 496 5076 504
rect 5148 496 5156 504
rect 5404 496 5412 504
rect 5500 496 5508 504
rect 5564 496 5572 504
rect 5772 496 5780 504
rect 5836 496 5844 504
rect 6220 496 6228 504
rect 1420 476 1428 484
rect 1660 476 1668 484
rect 1724 476 1732 484
rect 1932 476 1940 484
rect 1980 476 1988 484
rect 2508 476 2516 484
rect 3148 476 3156 484
rect 3180 476 3188 484
rect 3980 476 3988 484
rect 4044 476 4052 484
rect 4188 476 4196 484
rect 4332 476 4340 484
rect 4460 476 4468 484
rect 4476 476 4484 484
rect 4764 476 4772 484
rect 5180 476 5188 484
rect 5532 476 5540 484
rect 5580 476 5588 484
rect 5596 476 5604 484
rect 5612 476 5620 484
rect 6108 476 6116 484
rect 6204 476 6212 484
rect 300 456 308 464
rect 1004 456 1012 464
rect 1068 456 1076 464
rect 2524 456 2532 464
rect 3164 456 3172 464
rect 220 436 228 444
rect 460 436 468 444
rect 620 436 628 444
rect 924 436 932 444
rect 2940 436 2948 444
rect 3996 436 4004 444
rect 4028 436 4036 444
rect 4140 436 4148 444
rect 5164 436 5172 444
rect 5260 436 5268 444
rect 5436 436 5444 444
rect 5708 436 5716 444
rect 6156 436 6164 444
rect 1566 406 1574 414
rect 1580 406 1588 414
rect 1594 406 1602 414
rect 4638 406 4646 414
rect 4652 406 4660 414
rect 4666 406 4674 414
rect 492 376 500 384
rect 764 376 772 384
rect 796 376 804 384
rect 844 376 852 384
rect 1132 376 1140 384
rect 1324 376 1332 384
rect 1468 376 1476 384
rect 1532 376 1540 384
rect 1644 376 1652 384
rect 1692 376 1700 384
rect 1932 376 1940 384
rect 2028 376 2036 384
rect 2124 376 2132 384
rect 2892 376 2900 384
rect 2956 376 2964 384
rect 3356 376 3364 384
rect 3692 376 3700 384
rect 3884 376 3892 384
rect 4284 376 4292 384
rect 4364 376 4372 384
rect 4540 376 4548 384
rect 5100 376 5108 384
rect 5868 376 5876 384
rect 6044 376 6052 384
rect 6236 376 6244 384
rect 44 356 52 364
rect 556 356 564 364
rect 1196 356 1204 364
rect 1884 356 1892 364
rect 2588 356 2596 364
rect 3948 356 3956 364
rect 4124 356 4132 364
rect 6204 356 6212 364
rect 60 336 68 344
rect 236 336 244 344
rect 348 336 356 344
rect 476 336 484 344
rect 540 336 548 344
rect 1068 336 1076 344
rect 1084 336 1092 344
rect 1116 336 1124 344
rect 1180 336 1188 344
rect 1260 336 1268 344
rect 1308 336 1316 344
rect 1372 336 1380 344
rect 60 316 68 324
rect 204 316 212 324
rect 380 316 388 324
rect 508 316 516 324
rect 572 316 580 324
rect 732 316 740 324
rect 828 316 836 324
rect 956 316 964 324
rect 1020 316 1028 324
rect 1036 316 1044 324
rect 1148 316 1156 324
rect 1212 316 1220 324
rect 1228 316 1236 324
rect 1340 316 1348 324
rect 1436 336 1444 344
rect 1452 336 1460 344
rect 1516 336 1524 344
rect 1628 336 1636 344
rect 1676 336 1684 344
rect 1836 336 1844 344
rect 2716 336 2724 344
rect 3420 336 3428 344
rect 3932 336 3940 344
rect 4348 336 4356 344
rect 5404 336 5412 344
rect 5548 336 5556 344
rect 5916 336 5924 344
rect 1420 316 1428 324
rect 1484 316 1492 324
rect 1596 316 1604 324
rect 1708 316 1716 324
rect 1740 316 1748 324
rect 1788 316 1796 324
rect 1900 316 1908 324
rect 2140 316 2148 324
rect 2252 316 2260 324
rect 44 296 52 304
rect 76 296 84 304
rect 140 296 148 304
rect 220 296 228 304
rect 316 296 324 304
rect 364 296 372 304
rect 396 296 404 304
rect 492 296 500 304
rect 556 296 564 304
rect 636 296 644 304
rect 652 296 660 304
rect 796 296 804 304
rect 908 296 916 304
rect 972 296 980 304
rect 988 296 996 304
rect 1052 296 1060 304
rect 1132 296 1140 304
rect 1196 296 1204 304
rect 1244 296 1252 304
rect 1324 296 1332 304
rect 1388 296 1396 304
rect 1436 296 1444 304
rect 1500 296 1508 304
rect 1612 296 1620 304
rect 1692 296 1700 304
rect 1836 296 1844 304
rect 1932 296 1940 304
rect 2236 296 2244 304
rect 2428 316 2436 324
rect 2636 316 2644 324
rect 2764 316 2772 324
rect 2860 316 2868 324
rect 3212 316 3220 324
rect 3372 316 3380 324
rect 3580 316 3588 324
rect 3660 316 3668 324
rect 3836 316 3844 324
rect 3964 316 3972 324
rect 4044 316 4052 324
rect 4108 316 4116 324
rect 4316 316 4324 324
rect 4476 316 4484 324
rect 4572 316 4580 324
rect 4604 316 4612 324
rect 5132 316 5140 324
rect 5148 316 5156 324
rect 5180 316 5188 324
rect 5404 316 5412 324
rect 5452 316 5460 324
rect 5516 316 5524 324
rect 5580 316 5588 324
rect 5644 316 5652 324
rect 5820 316 5828 324
rect 5900 316 5908 324
rect 5996 316 6004 324
rect 6220 316 6228 324
rect 2460 296 2468 304
rect 2556 296 2564 304
rect 2652 296 2660 304
rect 2812 296 2820 304
rect 2892 296 2900 304
rect 3180 296 3188 304
rect 3596 296 3604 304
rect 3660 296 3668 304
rect 3692 296 3700 304
rect 3788 296 3796 304
rect 3868 296 3876 304
rect 3948 296 3956 304
rect 3980 296 3988 304
rect 4092 296 4100 304
rect 4140 296 4148 304
rect 92 276 100 284
rect 156 276 164 284
rect 300 276 308 284
rect 412 276 420 284
rect 620 276 628 284
rect 124 256 132 264
rect 188 256 196 264
rect 268 256 276 264
rect 364 256 372 264
rect 444 256 452 264
rect 588 256 596 264
rect 700 276 708 284
rect 780 276 788 284
rect 908 276 916 284
rect 972 276 980 284
rect 1276 276 1284 284
rect 1372 276 1380 284
rect 1852 276 1860 284
rect 1948 276 1956 284
rect 2060 276 2068 284
rect 2076 276 2084 284
rect 2108 276 2116 284
rect 2188 276 2196 284
rect 2364 276 2372 284
rect 2428 276 2436 284
rect 2460 276 2468 284
rect 2604 276 2612 284
rect 2652 276 2660 284
rect 2748 276 2756 284
rect 2796 276 2804 284
rect 2908 276 2916 284
rect 2924 276 2932 284
rect 3148 276 3156 284
rect 3228 276 3236 284
rect 3324 276 3332 284
rect 3340 276 3348 284
rect 3388 276 3396 284
rect 3484 276 3492 284
rect 3708 276 3716 284
rect 3804 276 3812 284
rect 3996 276 4004 284
rect 4028 276 4036 284
rect 4092 276 4100 284
rect 4140 276 4148 284
rect 4268 296 4276 304
rect 4364 296 4372 304
rect 4444 296 4452 304
rect 4460 296 4468 304
rect 4620 296 4628 304
rect 4780 296 4788 304
rect 4876 296 4884 304
rect 4940 296 4948 304
rect 5036 296 5044 304
rect 5068 296 5076 304
rect 5100 296 5108 304
rect 5196 296 5204 304
rect 5324 296 5332 304
rect 5340 296 5348 304
rect 5420 296 5428 304
rect 5500 296 5508 304
rect 5532 296 5540 304
rect 5612 296 5620 304
rect 5676 296 5684 304
rect 5756 296 5764 304
rect 5868 296 5876 304
rect 5916 296 5924 304
rect 6124 296 6132 304
rect 6172 296 6180 304
rect 4252 276 4260 284
rect 4268 276 4276 284
rect 748 256 756 264
rect 860 256 868 264
rect 876 256 884 264
rect 1724 256 1732 264
rect 1788 256 1796 264
rect 1868 256 1876 264
rect 2092 256 2100 264
rect 2156 256 2164 264
rect 2188 256 2196 264
rect 2284 256 2292 264
rect 2332 256 2340 264
rect 2476 256 2484 264
rect 2844 256 2852 264
rect 3036 256 3044 264
rect 3068 256 3076 264
rect 3500 256 3508 264
rect 3516 256 3524 264
rect 3532 256 3540 264
rect 3644 256 3652 264
rect 3740 256 3748 264
rect 3756 256 3764 264
rect 3900 256 3908 264
rect 4012 256 4020 264
rect 4268 256 4276 264
rect 4300 256 4308 264
rect 4428 276 4436 284
rect 4524 276 4532 284
rect 4748 276 4756 284
rect 4924 276 4932 284
rect 5052 276 5060 284
rect 5084 276 5092 284
rect 5244 276 5252 284
rect 5356 276 5364 284
rect 5580 276 5588 284
rect 5628 276 5636 284
rect 5660 276 5668 284
rect 5692 276 5700 284
rect 5740 276 5748 284
rect 5884 276 5892 284
rect 5964 276 5972 284
rect 6012 276 6020 284
rect 6108 276 6116 284
rect 6252 276 6260 284
rect 4492 256 4500 264
rect 4588 256 4596 264
rect 4908 256 4916 264
rect 4988 256 4996 264
rect 5004 256 5012 264
rect 5020 256 5028 264
rect 5228 256 5236 264
rect 5388 256 5396 264
rect 5468 256 5476 264
rect 5708 256 5716 264
rect 5932 256 5940 264
rect 5996 256 6004 264
rect 108 236 116 244
rect 172 236 180 244
rect 220 236 228 244
rect 284 236 292 244
rect 428 236 436 244
rect 604 236 612 244
rect 668 236 676 244
rect 1020 236 1028 244
rect 2764 236 2772 244
rect 2828 236 2836 244
rect 3292 236 3300 244
rect 3772 236 3780 244
rect 4636 236 4644 244
rect 4892 236 4900 244
rect 4972 236 4980 244
rect 5372 236 5380 244
rect 5484 236 5492 244
rect 5564 236 5572 244
rect 5740 236 5748 244
rect 6156 236 6164 244
rect 3118 206 3126 214
rect 3132 206 3140 214
rect 3146 206 3154 214
rect 204 176 212 184
rect 348 176 356 184
rect 860 176 868 184
rect 1004 176 1012 184
rect 1116 176 1124 184
rect 1276 176 1284 184
rect 1324 176 1332 184
rect 1388 176 1396 184
rect 1484 176 1492 184
rect 1804 176 1812 184
rect 1852 176 1860 184
rect 2300 176 2308 184
rect 2348 176 2356 184
rect 2476 176 2484 184
rect 2492 176 2500 184
rect 2764 176 2772 184
rect 2940 176 2948 184
rect 2988 176 2996 184
rect 3052 176 3060 184
rect 3516 176 3524 184
rect 3612 176 3620 184
rect 3676 176 3684 184
rect 4012 176 4020 184
rect 4156 176 4164 184
rect 4620 176 4628 184
rect 5132 176 5140 184
rect 5212 176 5220 184
rect 5436 176 5444 184
rect 5548 176 5556 184
rect 5948 176 5956 184
rect 6156 176 6164 184
rect 6204 176 6212 184
rect 332 156 340 164
rect 444 156 452 164
rect 460 156 468 164
rect 540 156 548 164
rect 556 156 564 164
rect 684 156 692 164
rect 956 156 964 164
rect 988 156 996 164
rect 1100 156 1108 164
rect 1292 156 1300 164
rect 1308 156 1316 164
rect 1404 156 1412 164
rect 1436 156 1444 164
rect 1500 156 1508 164
rect 1564 156 1572 164
rect 1916 156 1924 164
rect 1948 156 1956 164
rect 2028 156 2036 164
rect 2076 156 2084 164
rect 2220 156 2228 164
rect 2412 156 2420 164
rect 2604 156 2612 164
rect 2716 156 2724 164
rect 2748 156 2756 164
rect 2844 156 2852 164
rect 2924 156 2932 164
rect 2956 156 2964 164
rect 76 116 84 124
rect 140 136 148 144
rect 188 136 196 144
rect 252 136 260 144
rect 108 116 116 124
rect 236 116 244 124
rect 364 136 372 144
rect 508 136 516 144
rect 524 136 532 144
rect 652 136 660 144
rect 812 136 820 144
rect 988 136 996 144
rect 1020 136 1028 144
rect 1164 136 1172 144
rect 1260 136 1268 144
rect 1340 136 1348 144
rect 1436 136 1444 144
rect 1532 136 1540 144
rect 1628 136 1636 144
rect 1724 136 1732 144
rect 1740 136 1748 144
rect 1916 136 1924 144
rect 1980 136 1988 144
rect 2044 136 2052 144
rect 2188 136 2196 144
rect 2236 136 2244 144
rect 2332 136 2340 144
rect 2380 136 2388 144
rect 284 116 292 124
rect 380 116 388 124
rect 396 116 404 124
rect 492 116 500 124
rect 508 116 516 124
rect 588 116 596 124
rect 636 116 644 124
rect 732 116 740 124
rect 780 116 788 124
rect 796 116 804 124
rect 860 116 868 124
rect 908 116 916 124
rect 940 116 948 124
rect 1148 116 1156 124
rect 1244 116 1252 124
rect 1356 116 1364 124
rect 1452 116 1460 124
rect 2444 132 2452 140
rect 2588 136 2596 144
rect 2652 136 2660 144
rect 2700 136 2708 144
rect 2812 136 2820 144
rect 3196 156 3204 164
rect 3020 136 3028 144
rect 3052 136 3060 144
rect 3116 136 3124 144
rect 3308 156 3316 164
rect 3484 156 3492 164
rect 1884 116 1892 124
rect 1996 116 2004 124
rect 2012 116 2020 124
rect 2044 116 2052 124
rect 2188 116 2196 124
rect 2524 116 2532 124
rect 2620 116 2628 124
rect 2668 116 2676 124
rect 2716 116 2724 124
rect 2796 116 2804 124
rect 2892 116 2900 124
rect 2908 116 2916 124
rect 2972 116 2980 124
rect 3228 136 3236 144
rect 3452 136 3460 144
rect 3500 136 3508 144
rect 3548 136 3556 144
rect 3644 136 3652 144
rect 3692 136 3700 144
rect 3788 156 3796 164
rect 3868 156 3876 164
rect 3932 156 3940 164
rect 4076 156 4084 164
rect 4204 156 4212 164
rect 4300 156 4308 164
rect 4316 156 4324 164
rect 4364 156 4372 164
rect 4380 156 4388 164
rect 4428 156 4436 164
rect 4748 156 4756 164
rect 4844 156 4852 164
rect 4860 156 4868 164
rect 4924 156 4932 164
rect 5148 156 5156 164
rect 5196 156 5204 164
rect 5228 156 5236 164
rect 5308 156 5316 164
rect 5484 156 5492 164
rect 5644 156 5652 164
rect 5804 156 5812 164
rect 6220 156 6228 164
rect 3756 136 3764 144
rect 3788 136 3796 144
rect 3852 136 3860 144
rect 4044 136 4052 144
rect 4268 136 4276 144
rect 4364 136 4372 144
rect 4460 136 4468 144
rect 4780 136 4788 144
rect 4972 136 4980 144
rect 4988 136 4996 144
rect 5052 136 5060 144
rect 5084 136 5092 144
rect 5260 136 5268 144
rect 5388 136 5396 144
rect 5500 136 5508 144
rect 5548 136 5556 144
rect 5676 136 5684 144
rect 5708 136 5716 144
rect 5916 136 5924 144
rect 5932 136 5940 144
rect 5996 136 6004 144
rect 6172 136 6180 144
rect 3180 116 3188 124
rect 3212 116 3220 124
rect 3308 116 3316 124
rect 3340 116 3348 124
rect 3452 116 3460 124
rect 3708 116 3716 124
rect 3740 116 3748 124
rect 44 98 52 106
rect 188 96 196 104
rect 204 96 212 104
rect 316 96 324 104
rect 572 96 580 104
rect 684 96 692 104
rect 748 96 756 104
rect 764 96 772 104
rect 876 96 884 104
rect 604 76 612 84
rect 620 76 628 84
rect 716 76 724 84
rect 844 76 852 84
rect 1116 96 1124 104
rect 1228 96 1236 104
rect 1388 96 1396 104
rect 1484 96 1492 104
rect 1852 96 1860 104
rect 1932 96 1940 104
rect 1948 96 1956 104
rect 2348 96 2356 104
rect 2652 96 2660 104
rect 2764 96 2772 104
rect 2876 96 2884 104
rect 3052 96 3060 104
rect 3068 96 3076 104
rect 3260 96 3268 104
rect 3532 96 3540 104
rect 3660 96 3668 104
rect 3788 96 3796 104
rect 3836 116 3844 124
rect 4252 116 4260 124
rect 4284 96 4292 104
rect 4476 116 4484 124
rect 4524 116 4532 124
rect 4748 118 4756 126
rect 4812 116 4820 124
rect 4828 116 4836 124
rect 4892 116 4900 124
rect 5004 116 5012 124
rect 5068 116 5076 124
rect 5228 116 5236 124
rect 5340 116 5348 124
rect 5388 116 5396 124
rect 5436 116 5444 124
rect 5468 116 5476 124
rect 5564 116 5572 124
rect 5612 116 5620 124
rect 5660 116 5668 124
rect 5772 116 5780 124
rect 5932 116 5940 124
rect 6028 118 6036 126
rect 6172 116 6180 124
rect 4972 96 4980 104
rect 5036 96 5044 104
rect 5084 96 5092 104
rect 5308 96 5316 104
rect 5340 96 5348 104
rect 5452 96 5460 104
rect 5628 96 5636 104
rect 5964 96 5972 104
rect 924 76 932 84
rect 1068 76 1076 84
rect 4428 76 4436 84
rect 5372 76 5380 84
rect 5420 76 5428 84
rect 5596 76 5604 84
rect 284 56 292 64
rect 732 56 740 64
rect 5612 56 5620 64
rect 4508 36 4516 44
rect 4556 36 4564 44
rect 1566 6 1574 14
rect 1580 6 1588 14
rect 1594 6 1602 14
rect 4638 6 4646 14
rect 4652 6 4660 14
rect 4666 6 4674 14
<< metal2 >>
rect 237 5837 243 5843
rect 269 5837 275 5843
rect 493 5804 499 5843
rect 509 5837 531 5843
rect 781 5837 787 5843
rect 29 5684 35 5716
rect 45 5704 51 5716
rect 61 5704 67 5756
rect 157 5744 163 5756
rect 285 5744 291 5756
rect 301 5744 307 5756
rect 93 5703 99 5736
rect 84 5697 99 5703
rect 45 5564 51 5636
rect 77 5584 83 5696
rect 141 5584 147 5716
rect 221 5704 227 5736
rect 253 5724 259 5736
rect 189 5604 195 5676
rect 205 5584 211 5636
rect 237 5604 243 5716
rect 461 5704 467 5796
rect 509 5764 515 5837
rect 493 5704 499 5756
rect 509 5724 515 5756
rect 653 5744 659 5756
rect 669 5744 675 5776
rect 781 5724 787 5736
rect 589 5704 595 5716
rect 797 5703 803 5736
rect 813 5724 819 5843
rect 877 5837 883 5843
rect 829 5704 835 5796
rect 925 5764 931 5843
rect 845 5704 851 5716
rect 797 5697 812 5703
rect 285 5584 291 5596
rect 349 5544 355 5696
rect 605 5684 611 5696
rect 29 5517 44 5523
rect 29 5384 35 5517
rect 212 5517 220 5523
rect 61 5503 67 5516
rect 52 5497 67 5503
rect 13 5324 19 5376
rect 61 5244 67 5336
rect 77 5304 83 5496
rect 125 5384 131 5476
rect 141 5444 147 5496
rect 173 5484 179 5496
rect 189 5484 195 5496
rect 29 5184 35 5236
rect 93 5163 99 5316
rect 141 5184 147 5356
rect 157 5324 163 5336
rect 173 5324 179 5396
rect 205 5384 211 5456
rect 221 5364 227 5516
rect 237 5424 243 5496
rect 253 5464 259 5476
rect 93 5157 115 5163
rect 13 5064 19 5076
rect 61 4984 67 5096
rect 109 5043 115 5157
rect 221 5124 227 5276
rect 237 5244 243 5416
rect 253 5344 259 5456
rect 285 5444 291 5496
rect 269 5384 275 5436
rect 253 5184 259 5296
rect 285 5184 291 5336
rect 301 5324 307 5536
rect 717 5523 723 5556
rect 733 5544 739 5636
rect 717 5517 732 5523
rect 749 5504 755 5576
rect 477 5497 492 5503
rect 333 5464 339 5476
rect 349 5424 355 5496
rect 413 5444 419 5496
rect 445 5424 451 5456
rect 461 5444 467 5456
rect 349 5384 355 5396
rect 413 5357 451 5363
rect 413 5343 419 5357
rect 340 5337 355 5343
rect 212 5077 227 5083
rect 109 5037 131 5043
rect 125 4984 131 5037
rect 189 4984 195 5036
rect 221 4964 227 5077
rect 253 5044 259 5096
rect 269 5084 275 5116
rect 317 5083 323 5316
rect 349 5184 355 5337
rect 397 5337 419 5343
rect 397 5324 403 5337
rect 445 5324 451 5357
rect 477 5344 483 5497
rect 509 5464 515 5476
rect 621 5464 627 5476
rect 525 5344 531 5436
rect 541 5424 547 5436
rect 541 5344 547 5416
rect 589 5384 595 5436
rect 605 5364 611 5396
rect 765 5384 771 5536
rect 829 5404 835 5696
rect 868 5677 892 5683
rect 845 5664 851 5676
rect 845 5584 851 5656
rect 909 5644 915 5756
rect 925 5704 931 5756
rect 989 5744 995 5843
rect 1069 5804 1075 5843
rect 1133 5804 1139 5843
rect 1229 5837 1251 5843
rect 1021 5744 1027 5776
rect 1069 5744 1075 5796
rect 957 5704 963 5736
rect 909 5504 915 5536
rect 941 5523 947 5636
rect 989 5544 995 5736
rect 1021 5724 1027 5736
rect 1053 5724 1059 5736
rect 941 5517 963 5523
rect 957 5504 963 5517
rect 941 5464 947 5496
rect 1005 5484 1011 5716
rect 1021 5524 1027 5636
rect 1053 5604 1059 5696
rect 1085 5664 1091 5776
rect 1197 5744 1203 5756
rect 1133 5704 1139 5736
rect 1213 5704 1219 5756
rect 1101 5664 1107 5696
rect 1149 5644 1155 5696
rect 989 5424 995 5456
rect 1005 5444 1011 5476
rect 1005 5384 1011 5396
rect 845 5364 851 5376
rect 1069 5364 1075 5636
rect 1165 5604 1171 5636
rect 1101 5524 1107 5576
rect 1101 5404 1107 5496
rect 1133 5384 1139 5436
rect 1149 5384 1155 5436
rect 333 5104 339 5116
rect 381 5104 387 5116
rect 317 5077 339 5083
rect 333 4984 339 5077
rect 365 5064 371 5076
rect 381 5044 387 5076
rect 397 4984 403 5236
rect 413 5184 419 5316
rect 477 5304 483 5336
rect 493 5304 499 5336
rect 621 5324 627 5336
rect 452 5297 467 5303
rect 461 5104 467 5297
rect 493 5104 499 5296
rect 445 4984 451 5056
rect 461 4984 467 5096
rect 509 5064 515 5296
rect 541 5064 547 5316
rect 637 5184 643 5276
rect 717 5124 723 5356
rect 1133 5344 1139 5356
rect 829 5324 835 5336
rect 829 5184 835 5316
rect 925 5144 931 5336
rect 1037 5324 1043 5336
rect 1165 5304 1171 5596
rect 1213 5584 1219 5636
rect 1229 5524 1235 5837
rect 1293 5784 1299 5796
rect 1389 5764 1395 5843
rect 1453 5837 1475 5843
rect 1389 5744 1395 5756
rect 1325 5704 1331 5736
rect 1293 5584 1299 5616
rect 1325 5524 1331 5696
rect 1341 5624 1347 5736
rect 1405 5723 1411 5736
rect 1396 5717 1411 5723
rect 1357 5697 1372 5703
rect 1357 5604 1363 5697
rect 1421 5684 1427 5696
rect 1453 5684 1459 5837
rect 1501 5764 1507 5843
rect 1741 5837 1747 5843
rect 2077 5837 2083 5843
rect 2381 5837 2387 5843
rect 3037 5804 3043 5843
rect 3469 5837 3491 5843
rect 3112 5806 3118 5814
rect 3126 5806 3132 5814
rect 3140 5806 3146 5814
rect 3154 5806 3160 5814
rect 1469 5724 1475 5736
rect 1373 5604 1379 5656
rect 1293 5504 1299 5516
rect 1277 5484 1283 5496
rect 1261 5404 1267 5476
rect 1197 5344 1203 5356
rect 1053 5244 1059 5256
rect 893 5124 899 5136
rect 701 5084 707 5096
rect 541 4984 547 5056
rect 557 4984 563 5076
rect 76 4950 84 4956
rect 13 4684 19 4936
rect 77 4784 83 4796
rect 109 4684 115 4936
rect 157 4924 163 4936
rect 205 4924 211 4956
rect 221 4944 227 4956
rect 413 4944 419 4956
rect 573 4944 579 5036
rect 605 4984 611 5076
rect 765 5064 771 5116
rect 781 5064 787 5076
rect 893 5064 899 5076
rect 941 5064 947 5076
rect 893 4984 899 5056
rect 941 5024 947 5056
rect 957 4984 963 5096
rect 989 5084 995 5116
rect 1005 5084 1011 5096
rect 733 4944 739 4956
rect 925 4944 931 4976
rect 957 4964 963 4976
rect 317 4924 323 4936
rect 493 4924 499 4936
rect 173 4904 179 4916
rect 125 4804 131 4896
rect 13 4664 19 4676
rect 77 4584 83 4636
rect 109 4604 115 4676
rect 125 4583 131 4636
rect 125 4577 147 4583
rect 125 4544 131 4556
rect 13 4464 19 4536
rect 13 4284 19 4336
rect 45 4324 51 4376
rect 77 4184 83 4516
rect 109 4444 115 4536
rect 141 4524 147 4577
rect 189 4564 195 4656
rect 205 4543 211 4916
rect 381 4904 387 4916
rect 285 4884 291 4896
rect 493 4784 499 4916
rect 509 4904 515 4936
rect 669 4924 675 4936
rect 477 4704 483 4736
rect 637 4724 643 4736
rect 685 4724 691 4896
rect 717 4824 723 4936
rect 765 4884 771 4916
rect 893 4904 899 4916
rect 973 4903 979 4936
rect 973 4897 995 4903
rect 749 4784 755 4856
rect 237 4643 243 4676
rect 237 4637 259 4643
rect 221 4584 227 4596
rect 189 4537 211 4543
rect 157 4497 172 4503
rect 157 4304 163 4497
rect 141 4284 147 4296
rect 109 4264 115 4276
rect 189 4184 195 4537
rect 221 4384 227 4496
rect 237 4404 243 4536
rect 253 4184 259 4637
rect 349 4624 355 4676
rect 477 4664 483 4696
rect 269 4584 275 4616
rect 445 4584 451 4656
rect 493 4644 499 4696
rect 509 4664 515 4716
rect 525 4644 531 4716
rect 669 4684 675 4696
rect 685 4684 691 4716
rect 781 4684 787 4816
rect 893 4684 899 4716
rect 557 4664 563 4676
rect 621 4584 627 4616
rect 285 4524 291 4536
rect 269 4384 275 4496
rect 285 4483 291 4516
rect 285 4477 307 4483
rect 269 4244 275 4376
rect 285 4184 291 4456
rect 301 4264 307 4477
rect 397 4323 403 4536
rect 461 4504 467 4536
rect 461 4484 467 4496
rect 477 4464 483 4496
rect 493 4484 499 4576
rect 557 4504 563 4516
rect 573 4504 579 4556
rect 589 4484 595 4516
rect 605 4504 611 4536
rect 381 4317 403 4323
rect 317 4304 323 4316
rect 13 4124 19 4136
rect 125 4124 131 4136
rect 125 4083 131 4116
rect 125 4077 147 4083
rect 77 3984 83 4016
rect 125 3924 131 3936
rect 109 3884 115 3896
rect 13 3844 19 3876
rect 45 3784 51 3836
rect 125 3824 131 3916
rect 141 3904 147 4077
rect 189 3984 195 4056
rect 13 3704 19 3736
rect 77 3584 83 3716
rect 125 3704 131 3756
rect 157 3504 163 3896
rect 173 3784 179 3816
rect 205 3784 211 3896
rect 221 3804 227 4136
rect 269 4124 275 4136
rect 237 4084 243 4096
rect 285 4064 291 4096
rect 237 3904 243 3916
rect 260 3897 275 3903
rect 253 3884 259 3896
rect 269 3883 275 3897
rect 269 3877 284 3883
rect 237 3784 243 3836
rect 173 3584 179 3696
rect 164 3477 179 3483
rect 13 3344 19 3436
rect 45 3264 51 3296
rect 61 3184 67 3464
rect 109 3384 115 3476
rect 125 3384 131 3456
rect 173 3384 179 3477
rect 189 3384 195 3596
rect 221 3363 227 3516
rect 237 3384 243 3716
rect 253 3524 259 3856
rect 269 3724 275 3877
rect 285 3744 291 3856
rect 301 3744 307 4256
rect 269 3604 275 3716
rect 285 3604 291 3736
rect 317 3724 323 4276
rect 333 4144 339 4236
rect 381 4184 387 4317
rect 413 4303 419 4336
rect 429 4324 435 4356
rect 452 4337 467 4343
rect 413 4297 428 4303
rect 445 4284 451 4316
rect 461 4304 467 4337
rect 477 4284 483 4336
rect 573 4283 579 4336
rect 589 4324 595 4476
rect 605 4344 611 4496
rect 637 4384 643 4556
rect 653 4504 659 4636
rect 653 4484 659 4496
rect 589 4284 595 4316
rect 605 4304 611 4316
rect 564 4277 579 4283
rect 461 4184 467 4236
rect 493 4204 499 4236
rect 541 4164 547 4256
rect 333 4024 339 4116
rect 333 3724 339 3996
rect 349 3864 355 4136
rect 413 3904 419 3916
rect 413 3844 419 3876
rect 381 3784 387 3796
rect 413 3784 419 3816
rect 333 3704 339 3716
rect 301 3584 307 3636
rect 221 3357 243 3363
rect 173 3304 179 3356
rect 173 3224 179 3296
rect 205 3224 211 3336
rect 125 3124 131 3216
rect 221 3204 227 3296
rect 237 3184 243 3357
rect 253 3344 259 3516
rect 269 3504 275 3536
rect 333 3524 339 3596
rect 349 3584 355 3696
rect 365 3664 371 3716
rect 365 3584 371 3616
rect 333 3504 339 3516
rect 285 3364 291 3476
rect 333 3384 339 3496
rect 349 3384 355 3416
rect 365 3384 371 3556
rect 381 3464 387 3496
rect 397 3464 403 3596
rect 413 3584 419 3656
rect 429 3624 435 4036
rect 445 3984 451 4056
rect 493 4024 499 4136
rect 573 3984 579 4277
rect 637 4264 643 4296
rect 589 4184 595 4216
rect 637 4144 643 4256
rect 653 4164 659 4276
rect 589 4044 595 4116
rect 509 3864 515 3916
rect 493 3857 508 3863
rect 445 3644 451 3816
rect 461 3744 467 3756
rect 461 3704 467 3736
rect 477 3664 483 3696
rect 477 3604 483 3656
rect 493 3584 499 3857
rect 541 3824 547 3896
rect 589 3884 595 3956
rect 621 3924 627 4096
rect 669 3984 675 4656
rect 781 4644 787 4676
rect 877 4624 883 4656
rect 893 4604 899 4676
rect 829 4584 835 4596
rect 861 4544 867 4576
rect 973 4544 979 4576
rect 989 4564 995 4897
rect 1005 4744 1011 5056
rect 1037 4964 1043 5116
rect 1053 5104 1059 5236
rect 1069 5124 1075 5136
rect 1053 5064 1059 5076
rect 1101 5044 1107 5096
rect 1053 4984 1059 5036
rect 1085 4984 1091 4996
rect 1037 4924 1043 4956
rect 1069 4904 1075 4956
rect 1037 4884 1043 4896
rect 1085 4784 1091 4896
rect 1117 4804 1123 5076
rect 1133 5024 1139 5116
rect 1149 5104 1155 5296
rect 1181 5144 1187 5316
rect 1245 5304 1251 5376
rect 1181 5104 1187 5136
rect 1197 5124 1203 5296
rect 1245 5124 1251 5296
rect 1165 5044 1171 5096
rect 1181 5064 1187 5076
rect 1165 5004 1171 5036
rect 1197 4964 1203 5116
rect 1277 5084 1283 5456
rect 1293 5344 1299 5476
rect 1325 5444 1331 5516
rect 1341 5484 1347 5536
rect 1373 5524 1379 5596
rect 1405 5504 1411 5636
rect 1421 5504 1427 5576
rect 1453 5543 1459 5636
rect 1501 5604 1507 5756
rect 1517 5704 1523 5736
rect 1549 5704 1555 5796
rect 1844 5777 1987 5783
rect 1981 5764 1987 5777
rect 1517 5584 1523 5696
rect 1560 5606 1566 5614
rect 1574 5606 1580 5614
rect 1588 5606 1594 5614
rect 1602 5606 1608 5614
rect 1453 5537 1475 5543
rect 1437 5524 1443 5536
rect 1469 5524 1475 5537
rect 1389 5484 1395 5496
rect 1341 5464 1347 5476
rect 1389 5464 1395 5476
rect 1293 5284 1299 5336
rect 1357 5324 1363 5336
rect 1357 5123 1363 5316
rect 1405 5284 1411 5296
rect 1373 5184 1379 5276
rect 1437 5264 1443 5316
rect 1453 5304 1459 5516
rect 1581 5504 1587 5576
rect 1469 5424 1475 5436
rect 1469 5304 1475 5316
rect 1485 5304 1491 5316
rect 1501 5284 1507 5496
rect 1517 5344 1523 5476
rect 1533 5364 1539 5436
rect 1613 5364 1619 5496
rect 1629 5464 1635 5716
rect 1677 5704 1683 5756
rect 1725 5704 1731 5736
rect 1773 5724 1779 5756
rect 1821 5744 1827 5756
rect 1789 5624 1795 5696
rect 1805 5684 1811 5716
rect 1853 5624 1859 5756
rect 1965 5744 1971 5756
rect 1917 5737 1932 5743
rect 1869 5704 1875 5736
rect 1901 5704 1907 5736
rect 1917 5724 1923 5737
rect 1997 5724 2003 5756
rect 2004 5717 2019 5723
rect 1949 5684 1955 5716
rect 2013 5704 2019 5717
rect 2045 5703 2051 5716
rect 2077 5704 2083 5736
rect 2093 5724 2099 5736
rect 2141 5724 2147 5736
rect 2157 5724 2163 5756
rect 2205 5724 2211 5736
rect 2221 5724 2227 5756
rect 2029 5697 2051 5703
rect 2029 5684 2035 5697
rect 2125 5684 2131 5696
rect 2269 5684 2275 5696
rect 2285 5664 2291 5716
rect 2301 5684 2307 5716
rect 2349 5704 2355 5756
rect 2653 5744 2659 5756
rect 2717 5744 2723 5756
rect 3021 5744 3027 5756
rect 2381 5664 2387 5716
rect 1693 5484 1699 5516
rect 1885 5504 1891 5576
rect 1917 5504 1923 5616
rect 2157 5544 2163 5636
rect 1645 5424 1651 5456
rect 1709 5444 1715 5476
rect 1533 5344 1539 5356
rect 1565 5264 1571 5316
rect 1348 5117 1363 5123
rect 1325 5104 1331 5116
rect 1149 4904 1155 4916
rect 1165 4884 1171 4956
rect 1213 4924 1219 4996
rect 1229 4984 1235 5076
rect 1245 5024 1251 5036
rect 1245 5004 1251 5016
rect 1277 5004 1283 5076
rect 1309 5044 1315 5096
rect 1357 5064 1363 5076
rect 1373 5004 1379 5096
rect 1421 5064 1427 5076
rect 1421 5024 1427 5056
rect 1053 4664 1059 4696
rect 1085 4684 1091 4696
rect 1165 4684 1171 4696
rect 1005 4544 1011 4656
rect 1021 4584 1027 4636
rect 1037 4584 1043 4636
rect 1101 4584 1107 4596
rect 1133 4584 1139 4656
rect 1165 4624 1171 4656
rect 1181 4644 1187 4656
rect 1197 4644 1203 4676
rect 1229 4644 1235 4976
rect 1245 4944 1251 4956
rect 1437 4944 1443 5236
rect 1560 5206 1566 5214
rect 1574 5206 1580 5214
rect 1588 5206 1594 5214
rect 1602 5206 1608 5214
rect 1629 5104 1635 5416
rect 1645 5324 1651 5336
rect 1677 5283 1683 5436
rect 1725 5423 1731 5496
rect 1757 5484 1763 5496
rect 1773 5484 1779 5496
rect 1981 5484 1987 5536
rect 2045 5484 2051 5536
rect 1709 5417 1731 5423
rect 1668 5277 1683 5283
rect 1709 5264 1715 5417
rect 1725 5304 1731 5356
rect 1725 5224 1731 5296
rect 1741 5284 1747 5316
rect 1757 5284 1763 5436
rect 1693 5184 1699 5216
rect 1741 5104 1747 5116
rect 1757 5104 1763 5256
rect 1517 4944 1523 5036
rect 1597 4984 1603 5016
rect 1709 4984 1715 5036
rect 1492 4937 1507 4943
rect 1261 4924 1267 4936
rect 1309 4884 1315 4936
rect 1357 4904 1363 4936
rect 1405 4924 1411 4936
rect 1428 4897 1443 4903
rect 1293 4764 1299 4836
rect 1325 4804 1331 4836
rect 1373 4784 1379 4816
rect 1405 4784 1411 4836
rect 1293 4664 1299 4716
rect 1325 4704 1331 4736
rect 1389 4724 1395 4736
rect 1421 4704 1427 4736
rect 1437 4724 1443 4897
rect 1453 4824 1459 4916
rect 1453 4744 1459 4816
rect 1293 4624 1299 4656
rect 1341 4604 1347 4676
rect 1373 4664 1379 4696
rect 1405 4604 1411 4696
rect 1453 4684 1459 4696
rect 1469 4624 1475 4936
rect 1485 4884 1491 4916
rect 1501 4904 1507 4937
rect 1549 4904 1555 4936
rect 1581 4904 1587 4956
rect 1725 4944 1731 5056
rect 1773 4984 1779 5136
rect 1789 5064 1795 5436
rect 1837 5304 1843 5436
rect 1869 5424 1875 5476
rect 2125 5464 2131 5516
rect 2141 5504 2147 5536
rect 2205 5504 2211 5576
rect 2221 5544 2227 5636
rect 2285 5584 2291 5636
rect 2381 5544 2387 5636
rect 2285 5504 2291 5516
rect 2285 5484 2291 5496
rect 1901 5364 1907 5436
rect 1949 5384 1955 5456
rect 1997 5444 2003 5456
rect 2093 5384 2099 5396
rect 2221 5384 2227 5456
rect 2269 5364 2275 5436
rect 2301 5384 2307 5516
rect 2333 5484 2339 5536
rect 2413 5504 2419 5676
rect 2429 5644 2435 5736
rect 2541 5624 2547 5736
rect 2653 5704 2659 5736
rect 2749 5704 2755 5716
rect 2781 5704 2787 5716
rect 2573 5644 2579 5696
rect 2349 5464 2355 5476
rect 2317 5384 2323 5436
rect 2365 5364 2371 5496
rect 2445 5484 2451 5576
rect 2381 5464 2387 5476
rect 2429 5384 2435 5436
rect 1869 5324 1875 5336
rect 1917 5324 1923 5336
rect 1821 5264 1827 5296
rect 1853 5284 1859 5316
rect 1812 5077 1820 5083
rect 1789 5004 1795 5056
rect 1821 4944 1827 5076
rect 1837 5064 1843 5116
rect 1869 4944 1875 4976
rect 1901 4964 1907 5296
rect 1917 5143 1923 5276
rect 1965 5244 1971 5356
rect 2205 5324 2211 5336
rect 2125 5317 2140 5323
rect 1997 5244 2003 5296
rect 2013 5264 2019 5316
rect 2077 5184 2083 5276
rect 2093 5264 2099 5316
rect 2125 5184 2131 5317
rect 2189 5284 2195 5316
rect 2173 5184 2179 5256
rect 1917 5137 1939 5143
rect 1917 5084 1923 5096
rect 1917 4984 1923 4996
rect 1933 4984 1939 5137
rect 2141 5124 2147 5136
rect 2061 5104 2067 5116
rect 2189 5104 2195 5276
rect 2237 5244 2243 5356
rect 2397 5324 2403 5336
rect 2317 5304 2323 5316
rect 2253 5244 2259 5296
rect 2413 5284 2419 5356
rect 2445 5344 2451 5476
rect 2509 5424 2515 5436
rect 2541 5384 2547 5476
rect 2557 5464 2563 5636
rect 2573 5484 2579 5616
rect 2605 5584 2611 5676
rect 2813 5664 2819 5716
rect 2621 5644 2627 5656
rect 2861 5644 2867 5696
rect 2621 5484 2627 5636
rect 2653 5484 2659 5516
rect 2669 5484 2675 5496
rect 2701 5483 2707 5636
rect 2717 5524 2723 5636
rect 2877 5624 2883 5716
rect 2925 5684 2931 5736
rect 3133 5684 3139 5736
rect 3213 5704 3219 5736
rect 3229 5724 3235 5776
rect 3261 5724 3267 5736
rect 3357 5704 3363 5776
rect 3421 5724 3427 5776
rect 3469 5724 3475 5837
rect 3517 5744 3523 5843
rect 3821 5837 3843 5843
rect 3917 5837 3939 5843
rect 4029 5837 4035 5843
rect 4141 5837 4163 5843
rect 3837 5764 3843 5837
rect 3933 5764 3939 5837
rect 4141 5764 4147 5837
rect 3693 5724 3699 5756
rect 3213 5684 3219 5696
rect 3245 5684 3251 5696
rect 3389 5684 3395 5716
rect 3469 5704 3475 5716
rect 3405 5684 3411 5696
rect 2717 5484 2723 5516
rect 2749 5504 2755 5616
rect 2861 5544 2867 5556
rect 2909 5544 2915 5636
rect 3229 5544 3235 5636
rect 3245 5564 3251 5676
rect 2692 5477 2707 5483
rect 2733 5463 2739 5476
rect 2724 5457 2739 5463
rect 2477 5304 2483 5376
rect 2589 5364 2595 5456
rect 2621 5344 2627 5356
rect 2653 5304 2659 5316
rect 2685 5304 2691 5416
rect 2717 5364 2723 5456
rect 2749 5404 2755 5496
rect 2765 5324 2771 5496
rect 2829 5464 2835 5476
rect 2861 5444 2867 5496
rect 2941 5484 2947 5516
rect 3005 5504 3011 5536
rect 2797 5364 2803 5436
rect 2813 5364 2819 5376
rect 2845 5344 2851 5356
rect 2701 5304 2707 5316
rect 2781 5304 2787 5316
rect 2861 5304 2867 5316
rect 2877 5304 2883 5416
rect 2893 5324 2899 5356
rect 2909 5304 2915 5436
rect 2925 5424 2931 5456
rect 2957 5444 2963 5496
rect 3181 5484 3187 5496
rect 3213 5484 3219 5516
rect 3229 5504 3235 5536
rect 3277 5524 3283 5636
rect 3277 5504 3283 5516
rect 3293 5504 3299 5516
rect 3325 5484 3331 5636
rect 3437 5544 3443 5556
rect 3453 5544 3459 5636
rect 3341 5524 3347 5536
rect 3021 5444 3027 5476
rect 3053 5464 3059 5476
rect 2957 5324 2963 5356
rect 2669 5284 2675 5296
rect 2973 5284 2979 5436
rect 3069 5424 3075 5476
rect 3357 5464 3363 5496
rect 3421 5464 3427 5516
rect 3453 5504 3459 5536
rect 3437 5484 3443 5496
rect 3485 5484 3491 5516
rect 3112 5406 3118 5414
rect 3126 5406 3132 5414
rect 3140 5406 3146 5414
rect 3154 5406 3160 5414
rect 3181 5384 3187 5456
rect 3101 5344 3107 5356
rect 3197 5344 3203 5436
rect 3005 5324 3011 5336
rect 3021 5324 3027 5336
rect 3213 5324 3219 5376
rect 3325 5344 3331 5436
rect 3373 5384 3379 5436
rect 3341 5344 3347 5356
rect 2285 5124 2291 5236
rect 2493 5184 2499 5276
rect 2269 5117 2284 5123
rect 2205 5104 2211 5116
rect 2269 5084 2275 5117
rect 2093 5064 2099 5076
rect 2269 5064 2275 5076
rect 1933 4964 1939 4976
rect 1485 4704 1491 4796
rect 1501 4784 1507 4896
rect 1533 4764 1539 4896
rect 1629 4884 1635 4916
rect 1560 4806 1566 4814
rect 1574 4806 1580 4814
rect 1588 4806 1594 4814
rect 1602 4806 1608 4814
rect 1501 4737 1516 4743
rect 1501 4664 1507 4737
rect 1533 4684 1539 4696
rect 1501 4604 1507 4656
rect 1437 4584 1443 4596
rect 1517 4584 1523 4616
rect 1613 4584 1619 4756
rect 1629 4644 1635 4876
rect 1725 4844 1731 4936
rect 1821 4924 1827 4936
rect 1885 4924 1891 4936
rect 1853 4784 1859 4916
rect 1661 4684 1667 4736
rect 1677 4664 1683 4696
rect 1757 4684 1763 4736
rect 1773 4664 1779 4696
rect 1645 4624 1651 4656
rect 1597 4564 1603 4576
rect 685 4504 691 4516
rect 701 4504 707 4536
rect 717 4504 723 4516
rect 701 4384 707 4476
rect 685 4344 691 4356
rect 701 4304 707 4316
rect 717 4304 723 4316
rect 733 4184 739 4296
rect 749 4284 755 4316
rect 749 4184 755 4256
rect 765 4244 771 4496
rect 941 4484 947 4496
rect 989 4484 995 4516
rect 1005 4464 1011 4536
rect 1037 4504 1043 4556
rect 1069 4464 1075 4516
rect 829 4363 835 4396
rect 845 4384 851 4396
rect 829 4357 851 4363
rect 797 4304 803 4316
rect 813 4304 819 4316
rect 829 4264 835 4336
rect 813 4184 819 4236
rect 685 4104 691 4156
rect 749 4137 780 4143
rect 749 4123 755 4137
rect 740 4117 755 4123
rect 813 4104 819 4116
rect 829 4104 835 4256
rect 845 4244 851 4357
rect 909 4284 915 4436
rect 941 4264 947 4276
rect 845 4144 851 4236
rect 861 4144 867 4196
rect 877 4124 883 4216
rect 621 3803 627 3916
rect 669 3864 675 3916
rect 637 3824 643 3856
rect 621 3797 643 3803
rect 605 3784 611 3796
rect 637 3743 643 3797
rect 669 3784 675 3836
rect 685 3784 691 4096
rect 701 4084 707 4096
rect 701 4004 707 4076
rect 717 3984 723 4016
rect 797 3984 803 4036
rect 797 3904 803 3936
rect 813 3904 819 4096
rect 829 4044 835 4076
rect 829 3924 835 4036
rect 845 3984 851 4056
rect 701 3844 707 3896
rect 836 3877 851 3883
rect 813 3863 819 3876
rect 813 3857 835 3863
rect 749 3844 755 3856
rect 637 3737 659 3743
rect 525 3664 531 3696
rect 557 3644 563 3736
rect 573 3644 579 3736
rect 605 3684 611 3696
rect 429 3504 435 3516
rect 477 3504 483 3556
rect 557 3504 563 3556
rect 381 3424 387 3456
rect 397 3383 403 3456
rect 413 3424 419 3436
rect 429 3384 435 3456
rect 461 3424 467 3496
rect 477 3464 483 3496
rect 381 3377 403 3383
rect 253 3324 259 3336
rect 269 3284 275 3336
rect 173 3124 179 3176
rect 13 3044 19 3076
rect 164 3057 172 3063
rect 45 2944 51 3016
rect 93 2984 99 3036
rect 157 2944 163 3056
rect 173 2984 179 3036
rect 45 2784 51 2936
rect 93 2784 99 2816
rect 173 2764 179 2876
rect 189 2784 195 3036
rect 205 2984 211 3076
rect 253 3044 259 3076
rect 269 2984 275 3236
rect 285 3204 291 3336
rect 317 3304 323 3336
rect 349 3304 355 3336
rect 301 3264 307 3296
rect 365 3283 371 3296
rect 349 3277 371 3283
rect 285 3088 291 3196
rect 301 3163 307 3256
rect 317 3184 323 3256
rect 301 3157 323 3163
rect 285 2943 291 3080
rect 301 2944 307 2956
rect 276 2937 291 2943
rect 205 2884 211 2936
rect 221 2924 227 2936
rect 221 2824 227 2916
rect 237 2904 243 2936
rect 237 2784 243 2876
rect 269 2864 275 2936
rect 317 2924 323 3157
rect 333 3084 339 3216
rect 292 2917 307 2923
rect 109 2724 115 2736
rect 93 2584 99 2656
rect 109 2624 115 2716
rect 125 2543 131 2636
rect 173 2543 179 2756
rect 189 2544 195 2636
rect 205 2584 211 2676
rect 285 2644 291 2676
rect 301 2664 307 2917
rect 317 2904 323 2916
rect 333 2884 339 3076
rect 349 2984 355 3277
rect 381 3144 387 3377
rect 445 3364 451 3376
rect 413 3344 419 3356
rect 397 3264 403 3336
rect 397 3204 403 3256
rect 413 3183 419 3216
rect 445 3203 451 3356
rect 493 3344 499 3476
rect 525 3464 531 3476
rect 541 3464 547 3476
rect 477 3284 483 3336
rect 404 3177 419 3183
rect 429 3197 451 3203
rect 388 3097 403 3103
rect 397 3043 403 3097
rect 413 3064 419 3096
rect 397 3037 419 3043
rect 381 2984 387 3016
rect 413 2984 419 3037
rect 317 2704 323 2716
rect 349 2644 355 2956
rect 365 2824 371 2916
rect 429 2904 435 3197
rect 493 3144 499 3316
rect 525 3304 531 3416
rect 541 3344 547 3356
rect 509 3297 524 3303
rect 509 3104 515 3297
rect 541 3084 547 3336
rect 557 3324 563 3496
rect 573 3264 579 3556
rect 621 3524 627 3736
rect 653 3704 659 3737
rect 653 3663 659 3696
rect 653 3657 675 3663
rect 653 3504 659 3536
rect 669 3483 675 3657
rect 701 3584 707 3816
rect 749 3784 755 3836
rect 733 3724 739 3736
rect 765 3724 771 3796
rect 781 3744 787 3756
rect 797 3740 803 3796
rect 717 3564 723 3716
rect 653 3477 675 3483
rect 605 3404 611 3476
rect 621 3363 627 3456
rect 621 3357 643 3363
rect 605 3304 611 3316
rect 589 3284 595 3296
rect 477 3044 483 3076
rect 557 3063 563 3076
rect 541 3057 563 3063
rect 445 2924 451 2936
rect 477 2904 483 2916
rect 413 2864 419 2876
rect 397 2704 403 2776
rect 365 2684 371 2696
rect 365 2664 371 2676
rect 125 2537 147 2543
rect 13 2504 19 2516
rect 61 2504 67 2516
rect 109 2444 115 2496
rect 13 2184 19 2316
rect 45 2284 51 2436
rect 61 2324 67 2396
rect 93 2383 99 2436
rect 77 2377 99 2383
rect 45 2264 51 2276
rect 77 2263 83 2377
rect 93 2344 99 2356
rect 109 2284 115 2416
rect 125 2364 131 2516
rect 141 2484 147 2537
rect 157 2537 179 2543
rect 157 2463 163 2537
rect 173 2504 179 2516
rect 141 2457 163 2463
rect 141 2424 147 2457
rect 141 2284 147 2396
rect 157 2384 163 2436
rect 189 2404 195 2536
rect 237 2524 243 2636
rect 253 2584 259 2636
rect 269 2584 275 2636
rect 221 2504 227 2516
rect 269 2483 275 2576
rect 301 2524 307 2616
rect 349 2544 355 2556
rect 317 2504 323 2536
rect 269 2477 284 2483
rect 205 2364 211 2436
rect 157 2284 163 2356
rect 173 2317 188 2323
rect 157 2264 163 2276
rect 77 2257 99 2263
rect 29 2144 35 2236
rect 29 2084 35 2136
rect 45 2124 51 2236
rect 77 2224 83 2236
rect 93 2203 99 2257
rect 157 2244 163 2256
rect 77 2197 99 2203
rect 77 2104 83 2197
rect 109 2184 115 2236
rect 93 2124 99 2176
rect 109 2124 115 2176
rect 173 2164 179 2317
rect 221 2304 227 2476
rect 253 2364 259 2436
rect 301 2424 307 2436
rect 317 2344 323 2376
rect 333 2304 339 2416
rect 349 2344 355 2536
rect 381 2524 387 2636
rect 397 2464 403 2516
rect 349 2324 355 2336
rect 365 2304 371 2416
rect 237 2284 243 2296
rect 173 2144 179 2156
rect 13 1904 19 2036
rect 29 1884 35 1936
rect 61 1903 67 2096
rect 77 1924 83 2096
rect 93 1904 99 2116
rect 109 2084 115 2116
rect 61 1897 76 1903
rect 13 1704 19 1716
rect 45 1664 51 1836
rect 77 1764 83 1896
rect 93 1884 99 1896
rect 109 1863 115 2056
rect 125 1944 131 2036
rect 141 1904 147 1916
rect 157 1883 163 1896
rect 93 1857 115 1863
rect 141 1877 163 1883
rect 93 1784 99 1857
rect 61 1704 67 1716
rect 109 1704 115 1716
rect 45 1604 51 1636
rect 45 1484 51 1596
rect 13 1444 19 1476
rect 13 1364 19 1436
rect 45 924 51 936
rect 61 904 67 1576
rect 93 1504 99 1616
rect 125 1504 131 1836
rect 141 1804 147 1877
rect 141 1784 147 1796
rect 173 1744 179 1876
rect 189 1864 195 2216
rect 205 2204 211 2276
rect 253 2244 259 2276
rect 205 2140 211 2176
rect 205 1884 211 1956
rect 221 1944 227 2196
rect 253 2124 259 2196
rect 333 2164 339 2236
rect 269 1944 275 2136
rect 301 1944 307 1956
rect 333 1943 339 2036
rect 317 1937 339 1943
rect 221 1904 227 1936
rect 285 1904 291 1936
rect 189 1784 195 1836
rect 237 1724 243 1736
rect 157 1704 163 1716
rect 189 1644 195 1716
rect 253 1704 259 1816
rect 269 1724 275 1836
rect 269 1683 275 1716
rect 260 1677 275 1683
rect 189 1544 195 1636
rect 205 1504 211 1516
rect 77 924 83 1476
rect 93 1364 99 1496
rect 125 1484 131 1496
rect 141 1424 147 1436
rect 141 1323 147 1416
rect 132 1317 147 1323
rect 173 1284 179 1496
rect 237 1483 243 1636
rect 269 1624 275 1636
rect 269 1504 275 1556
rect 285 1484 291 1836
rect 301 1644 307 1756
rect 317 1503 323 1937
rect 333 1904 339 1916
rect 333 1724 339 1896
rect 349 1864 355 2296
rect 381 2284 387 2376
rect 413 2264 419 2336
rect 429 2304 435 2856
rect 493 2824 499 3056
rect 541 3004 547 3057
rect 541 2964 547 2996
rect 557 2984 563 3036
rect 573 3004 579 3256
rect 589 3044 595 3116
rect 605 3024 611 3276
rect 621 3064 627 3336
rect 637 3284 643 3357
rect 653 3344 659 3477
rect 701 3404 707 3456
rect 717 3424 723 3496
rect 733 3464 739 3716
rect 781 3684 787 3736
rect 813 3704 819 3796
rect 829 3784 835 3857
rect 845 3844 851 3877
rect 861 3824 867 4096
rect 893 4083 899 4156
rect 941 4124 947 4156
rect 957 4144 963 4196
rect 973 4124 979 4216
rect 893 4077 915 4083
rect 909 3984 915 4077
rect 877 3924 883 3936
rect 909 3924 915 3956
rect 941 3924 947 3936
rect 893 3884 899 3916
rect 909 3884 915 3896
rect 829 3737 844 3743
rect 829 3724 835 3737
rect 845 3704 851 3716
rect 861 3664 867 3776
rect 941 3704 947 3876
rect 957 3824 963 3876
rect 973 3804 979 3896
rect 957 3744 963 3756
rect 957 3704 963 3716
rect 797 3584 803 3656
rect 893 3644 899 3696
rect 957 3684 963 3696
rect 925 3584 931 3636
rect 765 3483 771 3516
rect 781 3504 787 3556
rect 829 3524 835 3536
rect 829 3504 835 3516
rect 765 3477 780 3483
rect 749 3424 755 3436
rect 669 3304 675 3396
rect 749 3384 755 3416
rect 685 3344 691 3356
rect 637 3043 643 3276
rect 653 3204 659 3296
rect 717 3284 723 3356
rect 653 3084 659 3156
rect 669 3122 675 3236
rect 733 3204 739 3316
rect 765 3284 771 3477
rect 797 3444 803 3496
rect 813 3444 819 3476
rect 829 3423 835 3496
rect 861 3484 867 3496
rect 893 3464 899 3576
rect 909 3524 915 3576
rect 813 3417 835 3423
rect 813 3384 819 3417
rect 781 3264 787 3336
rect 829 3324 835 3336
rect 788 3257 803 3263
rect 701 3104 707 3136
rect 797 3124 803 3257
rect 813 3204 819 3296
rect 829 3284 835 3316
rect 845 3224 851 3456
rect 973 3443 979 3576
rect 989 3464 995 4356
rect 1005 4304 1011 4336
rect 1021 4317 1036 4323
rect 1005 4184 1011 4296
rect 1021 4284 1027 4317
rect 1021 4184 1027 4276
rect 1053 4244 1059 4316
rect 1101 4264 1107 4556
rect 1117 4344 1123 4556
rect 1149 4483 1155 4536
rect 1165 4524 1171 4556
rect 1261 4544 1267 4556
rect 1133 4477 1155 4483
rect 1133 4324 1139 4477
rect 1165 4343 1171 4516
rect 1197 4403 1203 4536
rect 1188 4397 1203 4403
rect 1156 4337 1171 4343
rect 1037 4044 1043 4216
rect 1053 4204 1059 4236
rect 1069 4184 1075 4236
rect 1149 4184 1155 4336
rect 1181 4324 1187 4396
rect 1229 4384 1235 4516
rect 1309 4384 1315 4476
rect 1325 4444 1331 4516
rect 1341 4504 1347 4536
rect 1469 4504 1475 4516
rect 1213 4344 1219 4376
rect 1165 4304 1171 4316
rect 1245 4304 1251 4316
rect 1261 4304 1267 4376
rect 1421 4364 1427 4496
rect 1469 4384 1475 4496
rect 1485 4384 1491 4536
rect 1533 4384 1539 4536
rect 1725 4524 1731 4576
rect 1661 4444 1667 4516
rect 1741 4484 1747 4556
rect 1757 4504 1763 4536
rect 1560 4406 1566 4414
rect 1574 4406 1580 4414
rect 1588 4406 1594 4414
rect 1602 4406 1608 4414
rect 1165 4164 1171 4296
rect 1229 4284 1235 4296
rect 1277 4284 1283 4296
rect 1357 4284 1363 4316
rect 1309 4264 1315 4276
rect 1277 4144 1283 4176
rect 1053 4024 1059 4096
rect 1085 4064 1091 4136
rect 1069 3904 1075 3916
rect 1005 3704 1011 3776
rect 1021 3764 1027 3796
rect 1085 3784 1091 4036
rect 1101 4024 1107 4136
rect 1117 4064 1123 4116
rect 1101 3763 1107 3896
rect 1133 3884 1139 4136
rect 1213 4124 1219 4136
rect 1165 3924 1171 4116
rect 1181 4097 1196 4103
rect 1181 3924 1187 4097
rect 1229 4084 1235 4116
rect 1245 4104 1251 4116
rect 1309 4104 1315 4256
rect 1325 4224 1331 4276
rect 1421 4144 1427 4236
rect 1437 4204 1443 4316
rect 1485 4224 1491 4256
rect 1501 4184 1507 4276
rect 1549 4224 1555 4276
rect 1581 4204 1587 4316
rect 1645 4264 1651 4316
rect 1661 4304 1667 4316
rect 1709 4284 1715 4316
rect 1789 4304 1795 4756
rect 1901 4744 1907 4956
rect 1933 4944 1939 4956
rect 1981 4924 1987 4956
rect 1805 4624 1811 4716
rect 1869 4664 1875 4716
rect 1885 4704 1891 4736
rect 1901 4684 1907 4696
rect 1917 4684 1923 4896
rect 1933 4784 1939 4836
rect 1965 4744 1971 4916
rect 1981 4824 1987 4836
rect 1981 4784 1987 4796
rect 2013 4744 2019 4896
rect 2045 4864 2051 5056
rect 2061 4924 2067 4996
rect 2141 4944 2147 5016
rect 2173 4984 2179 5056
rect 2317 5044 2323 5096
rect 2365 5084 2371 5096
rect 2253 5024 2259 5036
rect 2189 4964 2195 5016
rect 2061 4784 2067 4876
rect 2077 4784 2083 4896
rect 2093 4884 2099 4936
rect 2141 4924 2147 4936
rect 2157 4924 2163 4936
rect 2125 4884 2131 4896
rect 2221 4884 2227 5016
rect 2285 4984 2291 5036
rect 2237 4924 2243 4936
rect 2253 4904 2259 4916
rect 2285 4884 2291 4976
rect 2301 4944 2307 4956
rect 2301 4924 2307 4936
rect 2317 4904 2323 4956
rect 2333 4924 2339 4976
rect 1965 4704 1971 4736
rect 1997 4724 2003 4736
rect 1981 4684 1987 4696
rect 1853 4544 1859 4556
rect 1869 4504 1875 4656
rect 1821 4384 1827 4436
rect 1901 4384 1907 4496
rect 1965 4444 1971 4556
rect 1997 4524 2003 4536
rect 1981 4504 1987 4516
rect 1981 4444 1987 4476
rect 1741 4284 1747 4296
rect 1869 4284 1875 4316
rect 1645 4184 1651 4256
rect 1853 4224 1859 4280
rect 1869 4264 1875 4276
rect 1917 4224 1923 4276
rect 1741 4184 1747 4196
rect 1949 4184 1955 4336
rect 1965 4304 1971 4356
rect 1981 4324 1987 4376
rect 1997 4304 2003 4356
rect 2013 4284 2019 4376
rect 2045 4344 2051 4736
rect 2077 4664 2083 4776
rect 2125 4744 2131 4796
rect 2141 4704 2147 4816
rect 2205 4724 2211 4876
rect 2301 4864 2307 4876
rect 2221 4684 2227 4696
rect 2141 4584 2147 4636
rect 2061 4484 2067 4536
rect 2109 4524 2115 4536
rect 2125 4524 2131 4536
rect 2077 4464 2083 4496
rect 2093 4484 2099 4496
rect 2157 4484 2163 4556
rect 2173 4544 2179 4556
rect 2189 4524 2195 4576
rect 2237 4503 2243 4556
rect 2228 4497 2243 4503
rect 2077 4344 2083 4356
rect 2093 4304 2099 4376
rect 1997 4184 2003 4256
rect 1565 4144 1571 4156
rect 1261 4084 1267 4096
rect 1236 4077 1251 4083
rect 1197 3984 1203 4056
rect 1165 3884 1171 3916
rect 1197 3904 1203 3956
rect 1245 3924 1251 4077
rect 1325 3984 1331 4096
rect 1277 3904 1283 3956
rect 1325 3884 1331 3896
rect 1117 3844 1123 3876
rect 1197 3844 1203 3876
rect 1213 3804 1219 3836
rect 1085 3757 1107 3763
rect 1021 3704 1027 3716
rect 973 3437 995 3443
rect 861 3384 867 3416
rect 861 3304 867 3356
rect 861 3164 867 3296
rect 893 3184 899 3396
rect 909 3304 915 3356
rect 941 3324 947 3416
rect 717 3084 723 3116
rect 861 3083 867 3116
rect 909 3103 915 3296
rect 909 3097 931 3103
rect 861 3077 876 3083
rect 653 3063 659 3076
rect 653 3057 675 3063
rect 621 3037 643 3043
rect 541 2943 547 2956
rect 525 2937 547 2943
rect 445 2724 451 2776
rect 509 2744 515 2836
rect 493 2664 499 2676
rect 445 2504 451 2636
rect 509 2624 515 2676
rect 461 2524 467 2536
rect 477 2504 483 2556
rect 509 2544 515 2556
rect 525 2543 531 2937
rect 541 2563 547 2716
rect 557 2684 563 2936
rect 573 2704 579 2996
rect 621 2984 627 3037
rect 589 2944 595 2976
rect 653 2964 659 3036
rect 605 2904 611 2916
rect 589 2684 595 2876
rect 637 2864 643 2936
rect 669 2924 675 3057
rect 685 2984 691 3076
rect 717 3044 723 3056
rect 717 2984 723 3036
rect 685 2844 691 2936
rect 749 2924 755 2996
rect 717 2884 723 2896
rect 637 2784 643 2816
rect 653 2763 659 2836
rect 701 2784 707 2836
rect 765 2804 771 3076
rect 861 3044 867 3077
rect 861 2984 867 3016
rect 781 2944 787 2956
rect 637 2757 659 2763
rect 612 2717 627 2723
rect 621 2684 627 2717
rect 557 2664 563 2676
rect 605 2624 611 2636
rect 541 2557 563 2563
rect 557 2544 563 2557
rect 525 2537 547 2543
rect 445 2484 451 2496
rect 445 2344 451 2476
rect 365 2104 371 2216
rect 381 2144 387 2216
rect 365 1884 371 1996
rect 397 1984 403 2236
rect 429 2163 435 2296
rect 445 2284 451 2316
rect 461 2304 467 2436
rect 429 2157 451 2163
rect 429 2004 435 2096
rect 445 1983 451 2157
rect 461 2123 467 2296
rect 477 2284 483 2336
rect 493 2304 499 2536
rect 509 2384 515 2496
rect 525 2444 531 2516
rect 541 2323 547 2537
rect 557 2504 563 2516
rect 573 2504 579 2536
rect 605 2524 611 2596
rect 621 2544 627 2656
rect 637 2564 643 2757
rect 653 2724 659 2736
rect 653 2604 659 2696
rect 669 2684 675 2756
rect 685 2704 691 2716
rect 621 2424 627 2536
rect 637 2344 643 2556
rect 669 2524 675 2536
rect 685 2524 691 2676
rect 701 2623 707 2776
rect 717 2744 723 2796
rect 797 2764 803 2936
rect 813 2864 819 2916
rect 829 2844 835 2936
rect 877 2923 883 3036
rect 909 2924 915 2936
rect 861 2917 883 2923
rect 765 2744 771 2756
rect 717 2724 723 2736
rect 749 2624 755 2736
rect 765 2704 771 2716
rect 765 2664 771 2696
rect 781 2664 787 2716
rect 797 2704 803 2716
rect 813 2624 819 2676
rect 829 2624 835 2636
rect 701 2617 723 2623
rect 717 2584 723 2617
rect 669 2364 675 2516
rect 669 2324 675 2356
rect 525 2317 547 2323
rect 477 2224 483 2236
rect 509 2204 515 2236
rect 477 2124 483 2136
rect 461 2117 476 2123
rect 493 2104 499 2156
rect 461 2084 467 2096
rect 461 2064 467 2076
rect 461 1984 467 1996
rect 429 1977 451 1983
rect 381 1884 387 1936
rect 365 1844 371 1876
rect 397 1784 403 1856
rect 349 1703 355 1736
rect 340 1697 355 1703
rect 349 1644 355 1676
rect 333 1564 339 1636
rect 365 1504 371 1716
rect 397 1564 403 1596
rect 429 1564 435 1977
rect 461 1964 467 1976
rect 477 1924 483 1936
rect 525 1904 531 2317
rect 557 2264 563 2276
rect 541 2124 547 2216
rect 589 2164 595 2276
rect 653 2264 659 2296
rect 557 2103 563 2136
rect 621 2124 627 2256
rect 605 2104 611 2116
rect 621 2104 627 2116
rect 637 2104 643 2156
rect 653 2124 659 2136
rect 541 2097 563 2103
rect 541 1984 547 2097
rect 477 1884 483 1896
rect 445 1784 451 1876
rect 461 1744 467 1756
rect 477 1740 483 1876
rect 445 1724 451 1736
rect 413 1504 419 1536
rect 477 1524 483 1676
rect 493 1644 499 1836
rect 509 1763 515 1836
rect 525 1824 531 1876
rect 509 1757 524 1763
rect 557 1744 563 1996
rect 573 1884 579 1916
rect 573 1764 579 1836
rect 509 1644 515 1716
rect 589 1704 595 1896
rect 621 1883 627 1996
rect 669 1943 675 2296
rect 685 2184 691 2316
rect 701 2304 707 2556
rect 749 2524 755 2536
rect 765 2524 771 2596
rect 813 2563 819 2596
rect 829 2584 835 2596
rect 813 2557 835 2563
rect 781 2504 787 2536
rect 813 2484 819 2536
rect 829 2524 835 2557
rect 845 2543 851 2736
rect 861 2724 867 2917
rect 861 2704 867 2716
rect 877 2604 883 2776
rect 893 2744 899 2896
rect 909 2864 915 2916
rect 925 2904 931 3097
rect 941 3064 947 3076
rect 957 2984 963 3316
rect 973 3184 979 3416
rect 989 3304 995 3437
rect 1005 3264 1011 3436
rect 1037 3384 1043 3496
rect 1069 3464 1075 3516
rect 1053 3424 1059 3456
rect 1085 3443 1091 3757
rect 1117 3724 1123 3776
rect 1133 3624 1139 3756
rect 1165 3704 1171 3716
rect 1197 3604 1203 3756
rect 1213 3744 1219 3796
rect 1357 3744 1363 4096
rect 1373 3884 1379 4136
rect 1405 4004 1411 4096
rect 1373 3864 1379 3876
rect 1405 3824 1411 3996
rect 1421 3984 1427 4136
rect 1444 4117 1459 4123
rect 1421 3864 1427 3916
rect 1453 3904 1459 4117
rect 1469 4064 1475 4096
rect 1581 4064 1587 4156
rect 1693 4144 1699 4156
rect 1709 4144 1715 4176
rect 1560 4006 1566 4014
rect 1574 4006 1580 4014
rect 1588 4006 1594 4014
rect 1602 4006 1608 4014
rect 1469 3884 1475 3936
rect 1133 3517 1148 3523
rect 1069 3437 1091 3443
rect 1037 3324 1043 3336
rect 1005 2984 1011 3056
rect 909 2744 915 2836
rect 925 2824 931 2876
rect 941 2844 947 2976
rect 932 2817 947 2823
rect 941 2704 947 2817
rect 893 2644 899 2676
rect 909 2664 915 2696
rect 957 2684 963 2856
rect 973 2704 979 2956
rect 989 2944 995 2956
rect 1021 2944 1027 3216
rect 1053 3204 1059 3276
rect 1037 3124 1043 3156
rect 1037 3104 1043 3116
rect 1053 3104 1059 3176
rect 1053 3084 1059 3096
rect 1021 2864 1027 2936
rect 1037 2924 1043 3056
rect 1069 2924 1075 3437
rect 1085 3304 1091 3316
rect 1101 3143 1107 3456
rect 1133 3404 1139 3517
rect 1181 3463 1187 3476
rect 1156 3457 1187 3463
rect 1149 3384 1155 3416
rect 1133 3144 1139 3156
rect 1101 3137 1123 3143
rect 1117 3123 1123 3137
rect 1165 3143 1171 3356
rect 1197 3324 1203 3596
rect 1245 3584 1251 3676
rect 1309 3644 1315 3736
rect 1373 3724 1379 3756
rect 1389 3724 1395 3736
rect 1277 3604 1283 3636
rect 1341 3584 1347 3716
rect 1373 3584 1379 3696
rect 1261 3544 1267 3556
rect 1229 3364 1235 3516
rect 1245 3504 1251 3536
rect 1277 3424 1283 3576
rect 1348 3557 1379 3563
rect 1293 3504 1299 3556
rect 1373 3544 1379 3557
rect 1309 3504 1315 3536
rect 1357 3504 1363 3516
rect 1389 3504 1395 3696
rect 1405 3524 1411 3796
rect 1421 3704 1427 3856
rect 1437 3764 1443 3836
rect 1485 3804 1491 3976
rect 1613 3884 1619 3896
rect 1629 3864 1635 4136
rect 1645 3984 1651 4096
rect 1661 3904 1667 4076
rect 1693 3984 1699 4136
rect 1805 4064 1811 4136
rect 1917 4124 1923 4156
rect 1949 4144 1955 4156
rect 1837 4084 1843 4116
rect 1869 4104 1875 4116
rect 1997 4104 2003 4116
rect 1837 4024 1843 4036
rect 1901 3924 1907 4036
rect 1997 4004 2003 4096
rect 1965 3984 1971 3996
rect 2013 3983 2019 4136
rect 2029 4004 2035 4216
rect 2045 4184 2051 4256
rect 2093 4224 2099 4236
rect 2109 4204 2115 4316
rect 2061 4124 2067 4136
rect 2109 4064 2115 4096
rect 2125 4044 2131 4156
rect 2004 3977 2019 3983
rect 2045 3904 2051 3916
rect 1613 3857 1628 3863
rect 1485 3744 1491 3796
rect 1437 3724 1443 3736
rect 1453 3703 1459 3716
rect 1501 3704 1507 3716
rect 1533 3704 1539 3716
rect 1581 3704 1587 3816
rect 1613 3704 1619 3857
rect 1709 3824 1715 3876
rect 1629 3784 1635 3816
rect 1709 3784 1715 3816
rect 1741 3744 1747 3836
rect 1773 3804 1779 3836
rect 1444 3697 1459 3703
rect 1421 3684 1427 3696
rect 1437 3644 1443 3676
rect 1469 3664 1475 3696
rect 1453 3523 1459 3636
rect 1560 3606 1566 3614
rect 1574 3606 1580 3614
rect 1588 3606 1594 3614
rect 1602 3606 1608 3614
rect 1533 3564 1539 3596
rect 1453 3517 1468 3523
rect 1421 3504 1427 3516
rect 1309 3484 1315 3496
rect 1341 3424 1347 3456
rect 1373 3424 1379 3496
rect 1421 3464 1427 3476
rect 1277 3384 1283 3396
rect 1309 3384 1315 3416
rect 1181 3284 1187 3316
rect 1181 3184 1187 3196
rect 1149 3137 1171 3143
rect 1117 3117 1139 3123
rect 1101 3083 1107 3116
rect 1092 3077 1107 3083
rect 1085 3064 1091 3076
rect 1069 2884 1075 2896
rect 1005 2744 1011 2836
rect 1037 2804 1043 2836
rect 1085 2764 1091 2956
rect 1133 2863 1139 3117
rect 1149 2984 1155 3137
rect 1165 3084 1171 3116
rect 1197 3004 1203 3236
rect 1229 3224 1235 3356
rect 1389 3344 1395 3396
rect 1437 3363 1443 3496
rect 1485 3484 1491 3496
rect 1501 3484 1507 3556
rect 1533 3464 1539 3556
rect 1565 3484 1571 3536
rect 1629 3524 1635 3696
rect 1645 3684 1651 3736
rect 1789 3724 1795 3816
rect 1805 3803 1811 3876
rect 1821 3864 1827 3896
rect 1869 3864 1875 3896
rect 1885 3864 1891 3876
rect 1821 3824 1827 3856
rect 1805 3797 1827 3803
rect 1757 3704 1763 3716
rect 1661 3584 1667 3656
rect 1645 3524 1651 3556
rect 1581 3484 1587 3516
rect 1469 3404 1475 3436
rect 1517 3384 1523 3396
rect 1421 3357 1443 3363
rect 1341 3324 1347 3336
rect 1373 3284 1379 3296
rect 1213 3024 1219 3116
rect 1229 3084 1235 3116
rect 1245 3104 1251 3236
rect 1165 2944 1171 2976
rect 1261 2924 1267 3236
rect 1277 3124 1283 3176
rect 1293 3043 1299 3236
rect 1325 3144 1331 3156
rect 1309 3104 1315 3136
rect 1341 3124 1347 3156
rect 1421 3144 1427 3357
rect 1453 3344 1459 3356
rect 1581 3264 1587 3416
rect 1597 3384 1603 3436
rect 1613 3424 1619 3496
rect 1661 3424 1667 3456
rect 1677 3384 1683 3696
rect 1805 3644 1811 3736
rect 1821 3724 1827 3797
rect 1837 3784 1843 3856
rect 1853 3844 1859 3856
rect 1981 3784 1987 3856
rect 1853 3764 1859 3776
rect 1885 3740 1891 3776
rect 1997 3764 2003 3896
rect 2077 3864 2083 4036
rect 2141 3944 2147 4336
rect 2189 4304 2195 4316
rect 2205 4284 2211 4456
rect 2237 4263 2243 4497
rect 2253 4444 2259 4636
rect 2269 4544 2275 4556
rect 2285 4524 2291 4576
rect 2269 4304 2275 4416
rect 2301 4324 2307 4636
rect 2317 4544 2323 4896
rect 2365 4844 2371 5076
rect 2413 5044 2419 5096
rect 2445 5084 2451 5096
rect 2429 5064 2435 5076
rect 2525 5024 2531 5116
rect 2573 5064 2579 5076
rect 2413 4884 2419 4996
rect 2429 4884 2435 4916
rect 2429 4764 2435 4836
rect 2461 4744 2467 4956
rect 2477 4884 2483 4996
rect 2493 4884 2499 4916
rect 2509 4904 2515 4976
rect 2541 4903 2547 5056
rect 2589 5044 2595 5096
rect 2557 4984 2563 5036
rect 2605 5004 2611 5076
rect 2621 5064 2627 5116
rect 2685 5044 2691 5096
rect 2733 5084 2739 5236
rect 2781 5083 2787 5236
rect 2893 5104 2899 5236
rect 2989 5104 2995 5236
rect 2980 5097 2988 5103
rect 2781 5077 2796 5083
rect 2557 4924 2563 4976
rect 2669 4964 2675 5036
rect 2701 4984 2707 5056
rect 2621 4924 2627 4956
rect 2733 4944 2739 4956
rect 2781 4944 2787 5036
rect 2861 4984 2867 5036
rect 2653 4924 2659 4936
rect 2797 4924 2803 4936
rect 2573 4904 2579 4916
rect 2589 4904 2595 4916
rect 2621 4904 2627 4916
rect 2532 4897 2547 4903
rect 2701 4884 2707 4896
rect 2717 4884 2723 4896
rect 2333 4584 2339 4696
rect 2333 4564 2339 4576
rect 2349 4504 2355 4656
rect 2365 4644 2371 4676
rect 2413 4564 2419 4636
rect 2397 4524 2403 4556
rect 2429 4544 2435 4656
rect 2413 4523 2419 4536
rect 2445 4524 2451 4636
rect 2461 4624 2467 4636
rect 2477 4603 2483 4716
rect 2493 4704 2499 4836
rect 2573 4724 2579 4756
rect 2621 4744 2627 4836
rect 2701 4744 2707 4776
rect 2628 4737 2636 4743
rect 2541 4684 2547 4716
rect 2573 4704 2579 4716
rect 2653 4704 2659 4716
rect 2669 4684 2675 4716
rect 2717 4704 2723 4876
rect 2813 4864 2819 4916
rect 2861 4903 2867 4956
rect 2925 4944 2931 4976
rect 2941 4944 2947 5036
rect 2861 4897 2876 4903
rect 2877 4884 2883 4896
rect 2461 4597 2483 4603
rect 2413 4517 2435 4523
rect 2429 4503 2435 4517
rect 2429 4497 2444 4503
rect 2260 4277 2275 4283
rect 2237 4257 2259 4263
rect 2205 4244 2211 4256
rect 2221 4204 2227 4256
rect 2212 4137 2227 4143
rect 2205 4084 2211 4116
rect 2221 4104 2227 4137
rect 2237 4124 2243 4136
rect 2253 4124 2259 4257
rect 2269 4244 2275 4277
rect 2157 3924 2163 4036
rect 2173 3903 2179 3916
rect 2189 3904 2195 4056
rect 2221 4024 2227 4096
rect 2269 4044 2275 4176
rect 2285 4163 2291 4316
rect 2349 4304 2355 4396
rect 2397 4384 2403 4436
rect 2461 4404 2467 4597
rect 2637 4584 2643 4656
rect 2669 4624 2675 4676
rect 2701 4584 2707 4616
rect 2621 4564 2627 4576
rect 2717 4563 2723 4636
rect 2717 4557 2739 4563
rect 2525 4504 2531 4536
rect 2589 4484 2595 4556
rect 2653 4524 2659 4536
rect 2669 4524 2675 4556
rect 2397 4324 2403 4336
rect 2429 4324 2435 4336
rect 2285 4157 2307 4163
rect 2301 4124 2307 4157
rect 2317 4144 2323 4276
rect 2333 4244 2339 4296
rect 2365 4284 2371 4316
rect 2445 4304 2451 4316
rect 2397 4284 2403 4296
rect 2413 4284 2419 4296
rect 2365 4144 2371 4216
rect 2397 4144 2403 4156
rect 2413 4144 2419 4156
rect 2445 4144 2451 4296
rect 2461 4104 2467 4196
rect 2477 4164 2483 4236
rect 2221 3984 2227 3996
rect 2205 3944 2211 3956
rect 2164 3897 2179 3903
rect 1933 3744 1939 3756
rect 1997 3744 2003 3756
rect 2061 3744 2067 3756
rect 1869 3724 1875 3736
rect 1981 3704 1987 3736
rect 2125 3704 2131 3796
rect 2173 3784 2179 3836
rect 2189 3744 2195 3796
rect 2237 3784 2243 3856
rect 2141 3724 2147 3736
rect 2189 3704 2195 3736
rect 1709 3604 1715 3636
rect 1693 3484 1699 3516
rect 1709 3504 1715 3596
rect 1693 3464 1699 3476
rect 1709 3464 1715 3496
rect 1741 3484 1747 3556
rect 1789 3544 1795 3596
rect 1805 3504 1811 3556
rect 1885 3504 1891 3636
rect 1933 3522 1939 3636
rect 1981 3584 1987 3696
rect 1965 3504 1971 3516
rect 1949 3463 1955 3476
rect 1949 3457 1964 3463
rect 1661 3323 1667 3336
rect 1677 3324 1683 3356
rect 1789 3344 1795 3456
rect 1853 3444 1859 3456
rect 1652 3317 1667 3323
rect 1773 3244 1779 3296
rect 1560 3206 1566 3214
rect 1574 3206 1580 3214
rect 1588 3206 1594 3214
rect 1602 3206 1608 3214
rect 1325 3104 1331 3116
rect 1277 3037 1299 3043
rect 1117 2857 1139 2863
rect 1005 2704 1011 2716
rect 845 2537 860 2543
rect 845 2523 851 2537
rect 836 2517 851 2523
rect 749 2464 755 2476
rect 845 2444 851 2496
rect 861 2484 867 2516
rect 893 2304 899 2596
rect 909 2464 915 2556
rect 925 2524 931 2636
rect 957 2524 963 2616
rect 973 2544 979 2636
rect 1021 2624 1027 2636
rect 1037 2523 1043 2756
rect 1101 2724 1107 2796
rect 1053 2704 1059 2716
rect 1069 2584 1075 2596
rect 1053 2544 1059 2556
rect 1037 2517 1059 2523
rect 925 2464 931 2496
rect 1037 2444 1043 2496
rect 957 2404 963 2436
rect 941 2304 947 2316
rect 765 2244 771 2256
rect 797 2244 803 2276
rect 749 2204 755 2236
rect 685 2164 691 2176
rect 765 2163 771 2236
rect 756 2157 771 2163
rect 701 2104 707 2116
rect 653 1937 675 1943
rect 637 1904 643 1916
rect 621 1877 636 1883
rect 477 1504 483 1516
rect 317 1497 332 1503
rect 237 1477 252 1483
rect 221 1464 227 1476
rect 205 1344 211 1456
rect 189 1317 204 1323
rect 109 1124 115 1276
rect 109 1104 115 1116
rect 93 1084 99 1096
rect 109 1064 115 1076
rect 93 964 99 1036
rect 125 984 131 1236
rect 157 984 163 1056
rect 109 924 115 936
rect 125 923 131 976
rect 116 917 131 923
rect 45 384 51 836
rect 61 724 67 896
rect 77 884 83 916
rect 84 877 92 883
rect 61 663 67 716
rect 61 657 76 663
rect 61 584 67 636
rect 93 584 99 636
rect 109 624 115 836
rect 141 724 147 896
rect 173 704 179 1256
rect 189 1124 195 1317
rect 221 1304 227 1376
rect 237 1364 243 1436
rect 237 1304 243 1336
rect 253 1324 259 1376
rect 301 1363 307 1436
rect 317 1384 323 1476
rect 301 1357 323 1363
rect 205 1124 211 1236
rect 237 1123 243 1296
rect 269 1284 275 1296
rect 301 1244 307 1336
rect 317 1324 323 1357
rect 333 1304 339 1496
rect 349 1424 355 1496
rect 365 1484 371 1496
rect 397 1484 403 1496
rect 509 1484 515 1496
rect 509 1464 515 1476
rect 349 1284 355 1296
rect 237 1117 252 1123
rect 269 1104 275 1116
rect 253 1097 268 1103
rect 189 1044 195 1056
rect 189 944 195 1036
rect 205 923 211 956
rect 196 917 211 923
rect 221 884 227 936
rect 237 924 243 936
rect 253 923 259 1097
rect 269 943 275 1076
rect 285 964 291 1036
rect 269 937 291 943
rect 253 917 275 923
rect 269 904 275 917
rect 253 884 259 896
rect 285 884 291 937
rect 301 924 307 1236
rect 349 1204 355 1276
rect 365 1264 371 1436
rect 397 1304 403 1316
rect 413 1304 419 1356
rect 445 1284 451 1436
rect 493 1404 499 1436
rect 525 1424 531 1696
rect 557 1504 563 1536
rect 541 1497 556 1503
rect 461 1304 467 1316
rect 477 1304 483 1336
rect 493 1304 499 1356
rect 525 1324 531 1396
rect 317 1084 323 1116
rect 365 1103 371 1236
rect 397 1104 403 1196
rect 461 1104 467 1236
rect 493 1184 499 1236
rect 509 1124 515 1316
rect 541 1144 547 1497
rect 573 1503 579 1636
rect 589 1624 595 1696
rect 573 1497 595 1503
rect 589 1444 595 1497
rect 605 1464 611 1756
rect 621 1584 627 1836
rect 637 1804 643 1876
rect 637 1724 643 1736
rect 653 1544 659 1937
rect 685 1904 691 2076
rect 717 2064 723 2136
rect 765 2084 771 2157
rect 813 2103 819 2276
rect 893 2263 899 2296
rect 916 2277 931 2283
rect 925 2264 931 2277
rect 884 2257 899 2263
rect 973 2263 979 2336
rect 1012 2317 1043 2323
rect 989 2304 995 2316
rect 1037 2304 1043 2317
rect 1037 2264 1043 2276
rect 948 2257 979 2263
rect 829 2124 835 2236
rect 861 2204 867 2236
rect 845 2144 851 2196
rect 877 2144 883 2176
rect 909 2124 915 2156
rect 925 2103 931 2256
rect 957 2184 963 2216
rect 813 2097 835 2103
rect 781 2064 787 2096
rect 733 1983 739 2036
rect 733 1977 755 1983
rect 749 1964 755 1977
rect 749 1904 755 1956
rect 813 1944 819 2036
rect 829 1984 835 2097
rect 909 2097 931 2103
rect 877 2004 883 2036
rect 909 1984 915 2097
rect 989 2064 995 2116
rect 1005 2104 1011 2156
rect 1037 2144 1043 2196
rect 1021 2124 1027 2136
rect 1053 2124 1059 2517
rect 1085 2504 1091 2716
rect 1101 2624 1107 2636
rect 1069 2384 1075 2436
rect 1069 2284 1075 2316
rect 1085 2244 1091 2296
rect 1117 2284 1123 2857
rect 1133 2804 1139 2836
rect 1133 2704 1139 2796
rect 1165 2704 1171 2716
rect 1181 2684 1187 2736
rect 1213 2684 1219 2696
rect 1149 2664 1155 2676
rect 1229 2664 1235 2676
rect 1165 2504 1171 2596
rect 1197 2583 1203 2636
rect 1245 2584 1251 2776
rect 1261 2704 1267 2796
rect 1277 2784 1283 3037
rect 1325 3024 1331 3096
rect 1341 2984 1347 3076
rect 1357 3064 1363 3096
rect 1373 3084 1379 3136
rect 1389 3064 1395 3136
rect 1421 3064 1427 3116
rect 1453 3104 1459 3156
rect 1469 3084 1475 3096
rect 1453 3064 1459 3076
rect 1501 3064 1507 3176
rect 1533 3144 1539 3176
rect 1549 3104 1555 3156
rect 1565 3104 1571 3116
rect 1629 3084 1635 3156
rect 1652 3137 1699 3143
rect 1661 3104 1667 3116
rect 1677 3064 1683 3116
rect 1693 3103 1699 3137
rect 1741 3104 1747 3236
rect 1805 3184 1811 3216
rect 1853 3164 1859 3436
rect 1869 3344 1875 3356
rect 1933 3344 1939 3396
rect 1869 3244 1875 3336
rect 1933 3304 1939 3336
rect 2013 3324 2019 3596
rect 2045 3584 2051 3656
rect 2173 3524 2179 3536
rect 2148 3517 2163 3523
rect 2052 3497 2076 3503
rect 2157 3424 2163 3517
rect 1773 3104 1779 3136
rect 1837 3124 1843 3136
rect 1869 3124 1875 3156
rect 1949 3144 1955 3236
rect 1965 3184 1971 3236
rect 1997 3164 2003 3236
rect 2013 3204 2019 3316
rect 2045 3124 2051 3296
rect 2077 3164 2083 3236
rect 2093 3144 2099 3316
rect 2157 3304 2163 3336
rect 2125 3264 2131 3296
rect 2173 3244 2179 3516
rect 2189 3504 2195 3536
rect 2205 3504 2211 3516
rect 2221 3484 2227 3496
rect 2237 3484 2243 3556
rect 2253 3463 2259 3876
rect 2269 3864 2275 3876
rect 2285 3823 2291 3896
rect 2301 3844 2307 3916
rect 2285 3817 2307 3823
rect 2269 3724 2275 3736
rect 2285 3724 2291 3756
rect 2301 3704 2307 3817
rect 2301 3584 2307 3696
rect 2317 3684 2323 4096
rect 2333 4044 2339 4096
rect 2461 4064 2467 4096
rect 2493 3884 2499 4436
rect 2509 4344 2515 4456
rect 2573 4364 2579 4436
rect 2653 4384 2659 4476
rect 2685 4424 2691 4556
rect 2733 4544 2739 4557
rect 2717 4464 2723 4536
rect 2717 4384 2723 4416
rect 2541 4264 2547 4296
rect 2557 4284 2563 4296
rect 2589 4264 2595 4336
rect 2733 4324 2739 4516
rect 2749 4464 2755 4696
rect 2765 4684 2771 4716
rect 2813 4684 2819 4856
rect 2845 4724 2851 4736
rect 2749 4384 2755 4436
rect 2765 4323 2771 4676
rect 2765 4317 2780 4323
rect 2605 4304 2611 4316
rect 2621 4264 2627 4296
rect 2509 4144 2515 4256
rect 2573 4204 2579 4236
rect 2356 3877 2371 3883
rect 2349 3724 2355 3756
rect 2365 3704 2371 3877
rect 2381 3804 2387 3856
rect 2397 3784 2403 3816
rect 2333 3684 2339 3696
rect 2349 3604 2355 3636
rect 2365 3624 2371 3696
rect 2381 3644 2387 3756
rect 2285 3504 2291 3536
rect 2301 3484 2307 3496
rect 2333 3464 2339 3496
rect 2349 3484 2355 3516
rect 2237 3457 2259 3463
rect 2237 3404 2243 3457
rect 2269 3444 2275 3456
rect 2189 3384 2195 3396
rect 2253 3344 2259 3436
rect 2317 3423 2323 3436
rect 2333 3424 2339 3456
rect 2301 3417 2323 3423
rect 2301 3384 2307 3417
rect 2317 3384 2323 3396
rect 2285 3324 2291 3336
rect 1693 3097 1708 3103
rect 1725 3064 1731 3076
rect 1389 3004 1395 3036
rect 1373 2944 1379 2976
rect 1389 2904 1395 2916
rect 1405 2904 1411 3056
rect 1517 3043 1523 3056
rect 1757 3044 1763 3076
rect 1501 3037 1523 3043
rect 1421 2924 1427 3036
rect 1485 3003 1491 3036
rect 1501 3003 1507 3037
rect 1485 2997 1507 3003
rect 1428 2917 1443 2923
rect 1325 2704 1331 2856
rect 1277 2697 1292 2703
rect 1277 2624 1283 2697
rect 1373 2684 1379 2696
rect 1293 2677 1308 2683
rect 1181 2577 1203 2583
rect 1133 2304 1139 2476
rect 1181 2424 1187 2577
rect 1277 2544 1283 2616
rect 1293 2544 1299 2677
rect 1389 2644 1395 2796
rect 1421 2784 1427 2836
rect 1405 2724 1411 2736
rect 1421 2684 1427 2736
rect 1437 2704 1443 2917
rect 1453 2904 1459 2956
rect 1485 2924 1491 2976
rect 1501 2944 1507 2997
rect 1517 2944 1523 2996
rect 1581 2944 1587 2996
rect 1613 2984 1619 2996
rect 1677 2984 1683 3016
rect 1693 2984 1699 3036
rect 1741 2944 1747 3036
rect 1789 2964 1795 3076
rect 1805 3064 1811 3096
rect 1853 3084 1859 3116
rect 1837 2984 1843 3056
rect 1869 3044 1875 3096
rect 1917 3044 1923 3096
rect 2045 3064 2051 3116
rect 2077 3104 2083 3116
rect 2093 3104 2099 3136
rect 2125 3083 2131 3156
rect 2189 3124 2195 3296
rect 2205 3284 2211 3296
rect 2205 3184 2211 3276
rect 2125 3077 2140 3083
rect 2237 3064 2243 3076
rect 1949 3057 1964 3063
rect 1533 2924 1539 2936
rect 1645 2924 1651 2936
rect 1805 2923 1811 2956
rect 1796 2917 1811 2923
rect 1620 2897 1628 2903
rect 1560 2806 1566 2814
rect 1574 2806 1580 2814
rect 1588 2806 1594 2814
rect 1602 2806 1608 2814
rect 1469 2724 1475 2736
rect 1341 2604 1347 2636
rect 1405 2624 1411 2636
rect 1389 2544 1395 2616
rect 1229 2484 1235 2496
rect 1069 2204 1075 2236
rect 1117 2184 1123 2276
rect 1181 2264 1187 2336
rect 1181 2144 1187 2236
rect 1197 2184 1203 2236
rect 1213 2164 1219 2176
rect 1229 2164 1235 2416
rect 1277 2324 1283 2516
rect 1405 2464 1411 2596
rect 1437 2524 1443 2576
rect 1437 2463 1443 2496
rect 1421 2457 1443 2463
rect 1245 2264 1251 2276
rect 1309 2264 1315 2316
rect 1037 2064 1043 2076
rect 1053 2063 1059 2116
rect 1181 2104 1187 2116
rect 1053 2057 1075 2063
rect 813 1904 819 1916
rect 692 1897 707 1903
rect 669 1784 675 1836
rect 685 1744 691 1816
rect 701 1764 707 1897
rect 733 1884 739 1896
rect 717 1804 723 1836
rect 717 1744 723 1776
rect 733 1743 739 1856
rect 765 1844 771 1876
rect 749 1764 755 1796
rect 733 1737 748 1743
rect 701 1724 707 1736
rect 669 1604 675 1716
rect 717 1644 723 1716
rect 733 1604 739 1716
rect 765 1704 771 1756
rect 781 1644 787 1836
rect 797 1764 803 1776
rect 813 1563 819 1836
rect 829 1684 835 1756
rect 845 1724 851 1816
rect 861 1684 867 1856
rect 893 1744 899 1916
rect 941 1904 947 2036
rect 1053 2004 1059 2036
rect 957 1924 963 1976
rect 1021 1884 1027 1996
rect 1069 1943 1075 2057
rect 1053 1937 1075 1943
rect 941 1864 947 1876
rect 909 1844 915 1856
rect 925 1824 931 1836
rect 941 1744 947 1756
rect 1021 1744 1027 1856
rect 1037 1804 1043 1916
rect 1053 1744 1059 1937
rect 1069 1824 1075 1836
rect 1069 1764 1075 1776
rect 925 1723 931 1736
rect 925 1717 940 1723
rect 877 1664 883 1716
rect 957 1704 963 1716
rect 797 1557 819 1563
rect 669 1504 675 1516
rect 797 1504 803 1557
rect 813 1524 819 1536
rect 621 1484 627 1496
rect 605 1424 611 1436
rect 557 1344 563 1396
rect 637 1384 643 1436
rect 653 1344 659 1496
rect 845 1484 851 1576
rect 861 1524 867 1636
rect 877 1584 883 1616
rect 893 1563 899 1656
rect 925 1584 931 1636
rect 989 1584 995 1736
rect 1085 1724 1091 2036
rect 1101 1944 1107 2016
rect 1117 1984 1123 2016
rect 1101 1924 1107 1936
rect 1133 1924 1139 1936
rect 1149 1904 1155 1996
rect 1213 1964 1219 2156
rect 1165 1884 1171 1936
rect 1117 1744 1123 1856
rect 1149 1744 1155 1856
rect 1005 1704 1011 1716
rect 877 1557 899 1563
rect 877 1504 883 1557
rect 893 1484 899 1536
rect 701 1464 707 1476
rect 717 1444 723 1480
rect 356 1097 371 1103
rect 365 1083 371 1097
rect 365 1077 380 1083
rect 333 944 339 976
rect 349 944 355 1036
rect 397 884 403 1096
rect 509 1084 515 1116
rect 541 1103 547 1136
rect 573 1124 579 1236
rect 621 1124 627 1156
rect 637 1104 643 1116
rect 653 1104 659 1336
rect 685 1304 691 1316
rect 701 1304 707 1316
rect 685 1244 691 1296
rect 733 1264 739 1456
rect 749 1364 755 1396
rect 765 1304 771 1456
rect 781 1364 787 1436
rect 829 1344 835 1416
rect 845 1324 851 1436
rect 781 1304 787 1316
rect 813 1304 819 1316
rect 541 1097 556 1103
rect 589 1084 595 1096
rect 653 1084 659 1096
rect 669 1084 675 1096
rect 685 1084 691 1196
rect 765 1184 771 1296
rect 701 1124 707 1156
rect 413 1064 419 1076
rect 429 1004 435 1036
rect 429 924 435 956
rect 493 924 499 956
rect 413 884 419 916
rect 477 884 483 916
rect 525 904 531 1036
rect 541 924 547 996
rect 605 884 611 1036
rect 621 924 627 996
rect 637 924 643 1036
rect 669 964 675 1036
rect 701 964 707 1036
rect 717 924 723 1176
rect 733 1104 739 1156
rect 749 1064 755 1076
rect 765 1043 771 1116
rect 797 1084 803 1176
rect 861 1164 867 1456
rect 877 1384 883 1396
rect 893 1364 899 1416
rect 909 1384 915 1536
rect 957 1484 963 1516
rect 925 1464 931 1476
rect 925 1404 931 1456
rect 925 1364 931 1376
rect 941 1304 947 1436
rect 973 1404 979 1576
rect 1005 1503 1011 1656
rect 1021 1524 1027 1676
rect 1037 1524 1043 1556
rect 1021 1504 1027 1516
rect 1069 1504 1075 1636
rect 1085 1544 1091 1716
rect 1101 1564 1107 1736
rect 1181 1724 1187 1956
rect 1229 1944 1235 1996
rect 1213 1924 1219 1936
rect 1197 1804 1203 1856
rect 1229 1804 1235 1896
rect 1245 1763 1251 2196
rect 1261 2124 1267 2236
rect 1277 2164 1283 2196
rect 1325 2123 1331 2416
rect 1421 2404 1427 2457
rect 1341 2304 1347 2336
rect 1437 2324 1443 2436
rect 1453 2424 1459 2616
rect 1469 2524 1475 2636
rect 1501 2624 1507 2796
rect 1533 2724 1539 2776
rect 1565 2704 1571 2776
rect 1517 2584 1523 2636
rect 1485 2544 1491 2576
rect 1453 2324 1459 2416
rect 1380 2317 1395 2323
rect 1364 2297 1379 2303
rect 1373 2244 1379 2297
rect 1389 2264 1395 2317
rect 1469 2303 1475 2376
rect 1485 2304 1491 2516
rect 1517 2484 1523 2556
rect 1533 2544 1539 2616
rect 1581 2584 1587 2676
rect 1629 2584 1635 2896
rect 1677 2864 1683 2896
rect 1709 2884 1715 2916
rect 1645 2724 1651 2756
rect 1693 2704 1699 2876
rect 1725 2864 1731 2916
rect 1741 2884 1747 2896
rect 1773 2884 1779 2916
rect 1789 2884 1795 2916
rect 1821 2903 1827 2956
rect 1853 2944 1859 2956
rect 1885 2924 1891 2996
rect 1933 2964 1939 2996
rect 1949 2984 1955 3057
rect 2045 3044 2051 3056
rect 1812 2897 1827 2903
rect 1837 2784 1843 2896
rect 1901 2844 1907 2936
rect 1949 2844 1955 2896
rect 1965 2884 1971 2996
rect 1997 2904 2003 3036
rect 2013 2924 2019 3016
rect 2061 2964 2067 2976
rect 2093 2884 2099 2976
rect 2109 2924 2115 3036
rect 2157 2984 2163 3036
rect 2205 3004 2211 3036
rect 2269 2984 2275 3256
rect 2317 3204 2323 3296
rect 2333 3224 2339 3416
rect 2365 3384 2371 3416
rect 2365 3324 2371 3356
rect 2349 3184 2355 3196
rect 2285 3064 2291 3116
rect 2397 3104 2403 3676
rect 2413 3664 2419 3736
rect 2461 3724 2467 3836
rect 2493 3784 2499 3876
rect 2509 3864 2515 4136
rect 2541 4124 2547 4176
rect 2557 4144 2563 4156
rect 2573 4104 2579 4156
rect 2637 4084 2643 4236
rect 2701 4184 2707 4256
rect 2701 4164 2707 4176
rect 2733 4144 2739 4196
rect 2653 4124 2659 4136
rect 2749 4124 2755 4176
rect 2541 3904 2547 3916
rect 2557 3884 2563 3936
rect 2605 3924 2611 3936
rect 2573 3884 2579 3916
rect 2509 3824 2515 3836
rect 2477 3744 2483 3756
rect 2573 3744 2579 3796
rect 2509 3724 2515 3736
rect 2573 3724 2579 3736
rect 2445 3704 2451 3716
rect 2429 3584 2435 3616
rect 2493 3524 2499 3676
rect 2413 3464 2419 3476
rect 2445 3464 2451 3496
rect 2477 3484 2483 3516
rect 2525 3504 2531 3636
rect 2557 3584 2563 3696
rect 2589 3684 2595 3836
rect 2605 3804 2611 3836
rect 2637 3784 2643 4036
rect 2653 3984 2659 4036
rect 2685 3984 2691 4096
rect 2653 3884 2659 3896
rect 2669 3804 2675 3876
rect 2701 3864 2707 4056
rect 2717 3924 2723 4036
rect 2749 3944 2755 4036
rect 2765 3944 2771 4276
rect 2797 4184 2803 4496
rect 2813 4464 2819 4496
rect 2829 4484 2835 4596
rect 2861 4524 2867 4756
rect 2909 4744 2915 4836
rect 2957 4744 2963 4996
rect 2973 4924 2979 5076
rect 3005 4983 3011 5316
rect 3181 5304 3187 5316
rect 3261 5284 3267 5336
rect 3357 5324 3363 5356
rect 3421 5324 3427 5336
rect 3277 5304 3283 5316
rect 3309 5304 3315 5316
rect 3293 5284 3299 5296
rect 3053 5124 3059 5136
rect 3149 5084 3155 5136
rect 3181 5103 3187 5236
rect 3245 5144 3251 5236
rect 3501 5184 3507 5276
rect 3309 5137 3324 5143
rect 3172 5097 3187 5103
rect 3165 5084 3171 5096
rect 3245 5084 3251 5116
rect 3053 5004 3059 5036
rect 3112 5006 3118 5014
rect 3126 5006 3132 5014
rect 3140 5006 3146 5014
rect 3154 5006 3160 5014
rect 2996 4977 3011 4983
rect 2989 4944 2995 4976
rect 3005 4944 3011 4956
rect 3181 4944 3187 4996
rect 3021 4764 3027 4836
rect 3037 4784 3043 4836
rect 3053 4763 3059 4896
rect 3197 4884 3203 5036
rect 3213 4984 3219 5076
rect 3293 5024 3299 5076
rect 3309 4984 3315 5137
rect 3325 5103 3331 5116
rect 3325 5097 3340 5103
rect 3325 5064 3331 5097
rect 3357 5024 3363 5116
rect 3373 4944 3379 4996
rect 3037 4757 3059 4763
rect 2957 4704 2963 4736
rect 2941 4684 2947 4696
rect 2957 4664 2963 4676
rect 2877 4544 2883 4596
rect 2813 4184 2819 4296
rect 2877 4284 2883 4396
rect 2893 4304 2899 4636
rect 2909 4484 2915 4556
rect 2813 4124 2819 4156
rect 2788 4117 2803 4123
rect 2797 4104 2803 4117
rect 2781 4064 2787 4096
rect 2813 3984 2819 4096
rect 2829 4084 2835 4196
rect 2861 4144 2867 4196
rect 2877 4084 2883 4236
rect 2893 4184 2899 4276
rect 2925 4264 2931 4536
rect 2941 4504 2947 4516
rect 2957 4424 2963 4536
rect 2973 4524 2979 4536
rect 2989 4504 2995 4716
rect 3005 4524 3011 4696
rect 3021 4664 3027 4736
rect 3005 4464 3011 4516
rect 3037 4423 3043 4757
rect 3053 4724 3059 4736
rect 3053 4544 3059 4656
rect 3069 4544 3075 4676
rect 3181 4664 3187 4856
rect 3112 4606 3118 4614
rect 3126 4606 3132 4614
rect 3140 4606 3146 4614
rect 3154 4606 3160 4614
rect 3181 4584 3187 4656
rect 3197 4564 3203 4876
rect 3213 4864 3219 4896
rect 3229 4884 3235 4916
rect 3389 4904 3395 5056
rect 3405 4944 3411 5116
rect 3421 5104 3427 5176
rect 3533 5164 3539 5436
rect 3581 5384 3587 5716
rect 3853 5704 3859 5756
rect 4061 5744 4067 5756
rect 4141 5744 4147 5756
rect 3885 5724 3891 5736
rect 4189 5724 4195 5843
rect 4253 5837 4259 5843
rect 4349 5837 4371 5843
rect 4365 5764 4371 5837
rect 4573 5837 4595 5843
rect 4573 5764 4579 5837
rect 4397 5724 4403 5756
rect 4685 5724 4691 5843
rect 5005 5837 5011 5843
rect 5037 5837 5043 5843
rect 5005 5764 5011 5776
rect 4749 5724 4755 5756
rect 3597 5484 3603 5576
rect 3741 5524 3747 5636
rect 3885 5584 3891 5636
rect 3645 5344 3651 5436
rect 3677 5324 3683 5496
rect 3773 5484 3779 5556
rect 3869 5484 3875 5496
rect 3885 5484 3891 5556
rect 3933 5524 3939 5716
rect 4093 5584 4099 5716
rect 4509 5704 4515 5716
rect 4605 5704 4611 5716
rect 4733 5684 4739 5716
rect 4765 5704 4771 5736
rect 4269 5584 4275 5656
rect 4285 5604 4291 5636
rect 4301 5524 4307 5536
rect 3933 5504 3939 5516
rect 3709 5477 3724 5483
rect 3709 5423 3715 5477
rect 3965 5463 3971 5516
rect 4109 5504 4115 5516
rect 4157 5504 4163 5516
rect 3997 5464 4003 5476
rect 3965 5457 3980 5463
rect 3693 5417 3715 5423
rect 3693 5344 3699 5417
rect 3517 5104 3523 5116
rect 3501 5084 3507 5096
rect 3421 5064 3427 5076
rect 3533 5064 3539 5136
rect 3549 5104 3555 5136
rect 3501 4984 3507 5036
rect 3533 4984 3539 5016
rect 3405 4924 3411 4936
rect 3229 4784 3235 4856
rect 3213 4644 3219 4736
rect 3261 4724 3267 4836
rect 3245 4704 3251 4716
rect 3229 4684 3235 4696
rect 3261 4684 3267 4696
rect 3261 4584 3267 4676
rect 3277 4644 3283 4676
rect 3229 4544 3235 4576
rect 3021 4417 3043 4423
rect 2717 3884 2723 3896
rect 2749 3884 2755 3916
rect 2765 3904 2771 3916
rect 2781 3904 2787 3916
rect 2589 3524 2595 3596
rect 2493 3384 2499 3476
rect 2525 3404 2531 3476
rect 2429 3324 2435 3356
rect 2445 3304 2451 3376
rect 2509 3304 2515 3376
rect 2541 3364 2547 3516
rect 2605 3483 2611 3636
rect 2621 3544 2627 3696
rect 2653 3584 2659 3616
rect 2701 3543 2707 3856
rect 2717 3784 2723 3836
rect 2765 3824 2771 3896
rect 2781 3784 2787 3856
rect 2765 3744 2771 3756
rect 2717 3737 2732 3743
rect 2717 3564 2723 3737
rect 2701 3537 2723 3543
rect 2605 3477 2620 3483
rect 2637 3404 2643 3476
rect 2573 3364 2579 3376
rect 2541 3324 2547 3336
rect 2653 3324 2659 3536
rect 2685 3504 2691 3516
rect 2701 3464 2707 3516
rect 2717 3463 2723 3537
rect 2733 3524 2739 3656
rect 2749 3624 2755 3716
rect 2765 3544 2771 3736
rect 2797 3644 2803 3936
rect 2829 3924 2835 4076
rect 2893 4044 2899 4096
rect 2813 3704 2819 3876
rect 2829 3844 2835 3876
rect 2829 3764 2835 3776
rect 2733 3484 2739 3516
rect 2765 3503 2771 3516
rect 2781 3504 2787 3516
rect 2756 3497 2771 3503
rect 2797 3464 2803 3536
rect 2829 3484 2835 3756
rect 2845 3744 2851 3796
rect 2877 3784 2883 3896
rect 2893 3844 2899 3876
rect 2893 3744 2899 3796
rect 2909 3784 2915 4256
rect 2925 4204 2931 4256
rect 2941 4144 2947 4236
rect 2957 4164 2963 4316
rect 2973 4304 2979 4336
rect 2957 4104 2963 4156
rect 2973 4124 2979 4196
rect 3021 4124 3027 4417
rect 3053 4384 3059 4496
rect 3085 4444 3091 4496
rect 3149 4484 3155 4536
rect 3277 4524 3283 4536
rect 3245 4504 3251 4516
rect 3181 4444 3187 4496
rect 3069 4424 3075 4436
rect 3197 4404 3203 4436
rect 3229 4384 3235 4436
rect 3261 4384 3267 4496
rect 3293 4484 3299 4716
rect 3309 4664 3315 4696
rect 3309 4484 3315 4656
rect 3325 4524 3331 4536
rect 3373 4504 3379 4796
rect 3389 4524 3395 4836
rect 3405 4804 3411 4876
rect 3421 4844 3427 4916
rect 3501 4864 3507 4896
rect 3469 4784 3475 4836
rect 3501 4784 3507 4816
rect 3405 4664 3411 4676
rect 3453 4664 3459 4736
rect 3501 4704 3507 4736
rect 3517 4683 3523 4896
rect 3533 4724 3539 4896
rect 3565 4784 3571 5036
rect 3581 4964 3587 5076
rect 3613 4964 3619 5156
rect 3629 5104 3635 5116
rect 3645 5104 3651 5116
rect 3661 5064 3667 5076
rect 3677 5064 3683 5296
rect 3693 5184 3699 5336
rect 3709 5144 3715 5316
rect 3725 5303 3731 5456
rect 3773 5324 3779 5336
rect 3757 5317 3772 5323
rect 3725 5297 3740 5303
rect 3741 5164 3747 5296
rect 3757 5184 3763 5317
rect 3805 5244 3811 5356
rect 3901 5324 3907 5416
rect 3821 5304 3827 5316
rect 3837 5284 3843 5316
rect 3853 5244 3859 5276
rect 3917 5204 3923 5436
rect 3949 5384 3955 5436
rect 3933 5363 3939 5376
rect 3933 5357 3948 5363
rect 3933 5304 3939 5357
rect 3869 5144 3875 5156
rect 3741 5104 3747 5136
rect 3693 5064 3699 5096
rect 3725 5084 3731 5096
rect 3677 4984 3683 5056
rect 3773 5044 3779 5096
rect 3789 5084 3795 5116
rect 3789 5064 3795 5076
rect 3821 4964 3827 5056
rect 3853 5044 3859 5136
rect 3933 5124 3939 5136
rect 3853 4984 3859 5016
rect 3869 4964 3875 5096
rect 3885 5044 3891 5116
rect 3613 4904 3619 4956
rect 3949 4944 3955 5196
rect 3965 5184 3971 5457
rect 4093 5444 4099 5476
rect 3997 5324 4003 5416
rect 4109 5384 4115 5496
rect 4157 5484 4163 5496
rect 4269 5444 4275 5496
rect 4333 5384 4339 5496
rect 4381 5464 4387 5536
rect 4093 5284 4099 5356
rect 4141 5324 4147 5356
rect 4109 5304 4115 5316
rect 4125 5304 4131 5316
rect 4157 5304 4163 5336
rect 4189 5324 4195 5356
rect 4205 5344 4211 5356
rect 4285 5304 4291 5336
rect 4317 5324 4323 5376
rect 4381 5324 4387 5436
rect 4397 5164 4403 5636
rect 4557 5584 4563 5676
rect 4632 5606 4638 5614
rect 4646 5606 4652 5614
rect 4660 5606 4666 5614
rect 4674 5606 4680 5614
rect 4733 5544 4739 5576
rect 4413 5344 4419 5516
rect 4477 5483 4483 5516
rect 4477 5477 4492 5483
rect 4429 5384 4435 5476
rect 4461 5344 4467 5356
rect 4461 5244 4467 5336
rect 4493 5304 4499 5476
rect 4525 5444 4531 5516
rect 4605 5504 4611 5516
rect 4525 5284 4531 5436
rect 4589 5384 4595 5476
rect 4605 5364 4611 5456
rect 4637 5444 4643 5516
rect 4701 5384 4707 5516
rect 4765 5484 4771 5696
rect 4861 5484 4867 5636
rect 4612 5357 4627 5363
rect 4573 5324 4579 5336
rect 4557 5304 4563 5316
rect 4621 5304 4627 5357
rect 4765 5356 4771 5476
rect 4877 5444 4883 5756
rect 4893 5704 4899 5756
rect 4925 5724 4931 5756
rect 4957 5664 4963 5716
rect 4973 5704 4979 5736
rect 5037 5724 5043 5776
rect 5357 5764 5363 5843
rect 5581 5764 5587 5843
rect 5149 5744 5155 5756
rect 5165 5724 5171 5736
rect 5053 5664 5059 5676
rect 4909 5524 4915 5556
rect 4781 5384 4787 5436
rect 4845 5344 4851 5436
rect 4925 5424 4931 5516
rect 4941 5504 4947 5536
rect 4957 5484 4963 5496
rect 5021 5484 5027 5536
rect 4989 5424 4995 5456
rect 4957 5384 4963 5416
rect 5053 5384 5059 5516
rect 5085 5503 5091 5636
rect 5133 5544 5139 5696
rect 5076 5497 5091 5503
rect 5117 5384 5123 5476
rect 4909 5344 4915 5376
rect 4701 5284 4707 5296
rect 4632 5206 4638 5214
rect 4646 5206 4652 5214
rect 4660 5206 4666 5214
rect 4674 5206 4680 5214
rect 4717 5184 4723 5256
rect 4797 5184 4803 5316
rect 4829 5184 4835 5316
rect 4845 5263 4851 5336
rect 4861 5304 4867 5336
rect 4909 5324 4915 5336
rect 4925 5324 4931 5356
rect 4973 5344 4979 5376
rect 5037 5324 5043 5356
rect 5053 5337 5068 5343
rect 4845 5257 4867 5263
rect 4061 5104 4067 5116
rect 3981 5044 3987 5076
rect 3789 4924 3795 4936
rect 3565 4704 3571 4736
rect 3597 4724 3603 4876
rect 3661 4844 3667 4916
rect 3709 4884 3715 4896
rect 3677 4864 3683 4876
rect 3725 4844 3731 4916
rect 3741 4864 3747 4876
rect 3773 4824 3779 4916
rect 3853 4824 3859 4936
rect 3885 4784 3891 4936
rect 3917 4904 3923 4936
rect 3949 4924 3955 4936
rect 3965 4924 3971 5036
rect 3997 5024 4003 5076
rect 4061 5064 4067 5096
rect 4045 5057 4060 5063
rect 3517 4677 3539 4683
rect 3037 4284 3043 4336
rect 3053 4304 3059 4316
rect 3085 4144 3091 4316
rect 3149 4284 3155 4336
rect 3181 4324 3187 4376
rect 3165 4304 3171 4316
rect 3181 4304 3187 4316
rect 3213 4284 3219 4336
rect 3277 4324 3283 4436
rect 3309 4384 3315 4456
rect 3357 4424 3363 4496
rect 3389 4484 3395 4496
rect 3405 4384 3411 4616
rect 3437 4584 3443 4636
rect 3469 4524 3475 4536
rect 3437 4483 3443 4496
rect 3428 4477 3443 4483
rect 3437 4424 3443 4477
rect 3229 4304 3235 4316
rect 3245 4244 3251 4316
rect 3112 4206 3118 4214
rect 3126 4206 3132 4214
rect 3140 4206 3146 4214
rect 3154 4206 3160 4214
rect 2925 3984 2931 4016
rect 2925 3844 2931 3856
rect 2941 3764 2947 4096
rect 2989 4064 2995 4076
rect 2973 3984 2979 4036
rect 2957 3924 2963 3936
rect 2877 3644 2883 3696
rect 2925 3604 2931 3696
rect 2941 3544 2947 3756
rect 2989 3683 2995 4056
rect 3005 3884 3011 3916
rect 3005 3864 3011 3876
rect 3021 3724 3027 4116
rect 3069 4044 3075 4096
rect 3085 4063 3091 4116
rect 3085 4057 3107 4063
rect 3037 3904 3043 3916
rect 3053 3904 3059 3916
rect 3101 3904 3107 4057
rect 3133 3984 3139 4176
rect 3181 4104 3187 4136
rect 3204 4117 3212 4123
rect 3245 4104 3251 4136
rect 3261 4083 3267 4296
rect 3277 4184 3283 4296
rect 3245 4077 3267 4083
rect 3245 3984 3251 4077
rect 3293 4063 3299 4336
rect 3357 4324 3363 4356
rect 3453 4344 3459 4496
rect 3469 4444 3475 4516
rect 3485 4423 3491 4496
rect 3469 4417 3491 4423
rect 3309 4184 3315 4196
rect 3309 4084 3315 4136
rect 3325 4124 3331 4276
rect 3357 4164 3363 4316
rect 3389 4304 3395 4336
rect 3405 4284 3411 4296
rect 3389 4277 3404 4283
rect 3389 4184 3395 4277
rect 3421 4144 3427 4236
rect 3469 4183 3475 4417
rect 3533 4244 3539 4677
rect 3549 4584 3555 4656
rect 3629 4604 3635 4736
rect 3789 4724 3795 4776
rect 3821 4724 3827 4736
rect 3645 4624 3651 4696
rect 3661 4664 3667 4716
rect 3773 4704 3779 4716
rect 3789 4704 3795 4716
rect 3677 4624 3683 4696
rect 3693 4604 3699 4676
rect 3549 4424 3555 4496
rect 3565 4384 3571 4596
rect 3741 4584 3747 4676
rect 3757 4663 3763 4696
rect 3757 4657 3772 4663
rect 3757 4564 3763 4576
rect 3821 4544 3827 4716
rect 3885 4664 3891 4716
rect 3933 4684 3939 4696
rect 3949 4684 3955 4696
rect 3933 4584 3939 4616
rect 3965 4584 3971 4896
rect 4013 4784 4019 4936
rect 4045 4904 4051 5057
rect 4093 4983 4099 5076
rect 4084 4977 4099 4983
rect 4077 4924 4083 4976
rect 4109 4963 4115 5096
rect 4141 4964 4147 5116
rect 4189 4984 4195 5156
rect 4221 5084 4227 5116
rect 4253 5064 4259 5136
rect 4461 5124 4467 5136
rect 4493 5124 4499 5176
rect 4525 5144 4531 5176
rect 4541 5124 4547 5156
rect 4573 5117 4643 5123
rect 4301 5104 4307 5116
rect 4100 4957 4115 4963
rect 4093 4944 4099 4956
rect 4221 4944 4227 5016
rect 4157 4904 4163 4936
rect 4205 4924 4211 4936
rect 4237 4924 4243 5036
rect 4285 4984 4291 5056
rect 4349 5044 4355 5076
rect 4397 5064 4403 5116
rect 4349 4984 4355 5036
rect 4269 4904 4275 4956
rect 4413 4924 4419 4936
rect 4061 4744 4067 4756
rect 4045 4604 4051 4736
rect 4077 4724 4083 4756
rect 4109 4684 4115 4696
rect 4141 4684 4147 4716
rect 4109 4584 4115 4616
rect 4141 4584 4147 4676
rect 4029 4544 4035 4556
rect 3581 4524 3587 4536
rect 3581 4384 3587 4516
rect 3533 4184 3539 4216
rect 3549 4184 3555 4336
rect 3565 4204 3571 4296
rect 3581 4264 3587 4316
rect 3572 4197 3587 4203
rect 3469 4177 3491 4183
rect 3485 4163 3491 4177
rect 3485 4157 3507 4163
rect 3277 4057 3299 4063
rect 3277 3984 3283 4057
rect 3325 4024 3331 4116
rect 3373 4084 3379 4136
rect 3389 4124 3395 4136
rect 3405 4064 3411 4096
rect 3421 4024 3427 4136
rect 3469 3944 3475 4096
rect 3485 3944 3491 3956
rect 3197 3904 3203 3916
rect 3277 3904 3283 3916
rect 3005 3684 3011 3696
rect 2989 3677 3004 3683
rect 2925 3484 2931 3536
rect 2973 3504 2979 3576
rect 2989 3504 2995 3556
rect 3005 3524 3011 3616
rect 3021 3524 3027 3716
rect 3037 3624 3043 3896
rect 3053 3804 3059 3896
rect 3085 3763 3091 3816
rect 3112 3806 3118 3814
rect 3126 3806 3132 3814
rect 3140 3806 3146 3814
rect 3154 3806 3160 3814
rect 3085 3757 3107 3763
rect 3069 3724 3075 3736
rect 3085 3724 3091 3736
rect 3085 3584 3091 3676
rect 3037 3544 3043 3556
rect 3053 3523 3059 3556
rect 3101 3544 3107 3757
rect 3181 3744 3187 3896
rect 3197 3824 3203 3876
rect 3245 3824 3251 3876
rect 3277 3824 3283 3896
rect 3309 3884 3315 3916
rect 3245 3784 3251 3816
rect 3309 3763 3315 3876
rect 3325 3784 3331 3876
rect 3341 3784 3347 3896
rect 3373 3824 3379 3916
rect 3357 3784 3363 3816
rect 3309 3757 3331 3763
rect 3181 3724 3187 3736
rect 3213 3724 3219 3756
rect 3117 3684 3123 3696
rect 3037 3517 3059 3523
rect 2973 3484 2979 3496
rect 3005 3484 3011 3516
rect 2941 3464 2947 3476
rect 2717 3457 2739 3463
rect 2717 3344 2723 3436
rect 2413 3204 2419 3276
rect 2429 3264 2435 3276
rect 2493 3264 2499 3296
rect 2525 3284 2531 3316
rect 2669 3284 2675 3296
rect 2189 2944 2195 2956
rect 2285 2944 2291 3056
rect 2301 2984 2307 3096
rect 2397 3084 2403 3096
rect 2317 3044 2323 3076
rect 2429 3063 2435 3116
rect 2461 3084 2467 3096
rect 2429 3057 2444 3063
rect 2317 2944 2323 3016
rect 2125 2904 2131 2936
rect 1741 2704 1747 2716
rect 1677 2684 1683 2696
rect 1661 2663 1667 2676
rect 1709 2663 1715 2696
rect 1757 2664 1763 2776
rect 1997 2744 2003 2836
rect 1789 2704 1795 2736
rect 1661 2657 1715 2663
rect 1741 2624 1747 2636
rect 1773 2564 1779 2636
rect 1789 2584 1795 2696
rect 1885 2684 1891 2716
rect 2029 2704 2035 2716
rect 1885 2664 1891 2676
rect 1901 2664 1907 2696
rect 1965 2684 1971 2696
rect 1981 2684 1987 2696
rect 1789 2544 1795 2576
rect 1805 2564 1811 2576
rect 1613 2524 1619 2536
rect 1661 2524 1667 2536
rect 1460 2297 1475 2303
rect 1501 2284 1507 2296
rect 1517 2284 1523 2316
rect 1533 2304 1539 2516
rect 1549 2484 1555 2516
rect 1693 2504 1699 2516
rect 1709 2504 1715 2536
rect 1805 2524 1811 2556
rect 1821 2544 1827 2636
rect 1869 2584 1875 2636
rect 1885 2504 1891 2596
rect 1901 2504 1907 2516
rect 1560 2406 1566 2414
rect 1574 2406 1580 2414
rect 1588 2406 1594 2414
rect 1602 2406 1608 2414
rect 1645 2304 1651 2396
rect 1565 2284 1571 2296
rect 1421 2244 1427 2276
rect 1517 2263 1523 2276
rect 1661 2264 1667 2436
rect 1677 2324 1683 2336
rect 1501 2257 1523 2263
rect 1357 2224 1363 2236
rect 1357 2143 1363 2216
rect 1405 2184 1411 2236
rect 1501 2204 1507 2257
rect 1517 2184 1523 2236
rect 1437 2144 1443 2176
rect 1357 2137 1379 2143
rect 1316 2117 1331 2123
rect 1277 2004 1283 2096
rect 1309 2084 1315 2096
rect 1341 2084 1347 2136
rect 1357 2084 1363 2116
rect 1373 2104 1379 2137
rect 1517 2104 1523 2156
rect 1533 2124 1539 2216
rect 1677 2164 1683 2236
rect 1629 2137 1667 2143
rect 1629 2124 1635 2137
rect 1661 2124 1667 2137
rect 1396 2097 1411 2103
rect 1293 1984 1299 2036
rect 1325 1924 1331 1936
rect 1325 1904 1331 1916
rect 1277 1864 1283 1876
rect 1229 1757 1251 1763
rect 1117 1717 1155 1723
rect 1117 1664 1123 1717
rect 1133 1664 1139 1696
rect 1149 1664 1155 1717
rect 1085 1504 1091 1536
rect 996 1497 1011 1503
rect 1069 1464 1075 1476
rect 1053 1424 1059 1436
rect 964 1377 979 1383
rect 973 1343 979 1377
rect 1021 1343 1027 1396
rect 1101 1384 1107 1496
rect 1133 1484 1139 1516
rect 1149 1484 1155 1636
rect 1165 1564 1171 1676
rect 1197 1604 1203 1696
rect 1181 1503 1187 1596
rect 1197 1524 1203 1536
rect 1172 1497 1187 1503
rect 973 1337 995 1343
rect 1021 1337 1036 1343
rect 957 1304 963 1336
rect 989 1324 995 1337
rect 1053 1304 1059 1356
rect 877 1284 883 1296
rect 861 1104 867 1156
rect 845 1084 851 1096
rect 749 1037 771 1043
rect 749 964 755 1037
rect 733 944 739 956
rect 749 944 755 956
rect 765 944 771 976
rect 781 944 787 1036
rect 797 984 803 1076
rect 861 1064 867 1076
rect 893 1043 899 1296
rect 909 1123 915 1196
rect 925 1143 931 1236
rect 941 1184 947 1236
rect 989 1224 995 1236
rect 973 1143 979 1176
rect 1069 1164 1075 1376
rect 1101 1323 1107 1376
rect 1092 1317 1107 1323
rect 1133 1264 1139 1476
rect 925 1137 947 1143
rect 973 1137 995 1143
rect 941 1124 947 1137
rect 909 1117 931 1123
rect 909 1084 915 1096
rect 925 1084 931 1117
rect 957 1097 972 1103
rect 957 1084 963 1097
rect 989 1084 995 1137
rect 989 1064 995 1076
rect 877 1037 899 1043
rect 813 964 819 1036
rect 845 964 851 976
rect 237 784 243 836
rect 285 704 291 836
rect 276 697 284 703
rect 205 684 211 696
rect 93 544 99 556
rect 109 544 115 556
rect 125 444 131 636
rect 221 624 227 676
rect 141 564 147 576
rect 189 504 195 536
rect 205 504 211 576
rect 221 524 227 616
rect 237 504 243 676
rect 253 604 259 636
rect 269 524 275 696
rect 301 683 307 776
rect 292 677 307 683
rect 301 524 307 677
rect 317 664 323 736
rect 333 724 339 776
rect 381 743 387 836
rect 429 744 435 836
rect 493 784 499 836
rect 541 744 547 836
rect 381 737 403 743
rect 397 704 403 737
rect 461 724 467 736
rect 397 664 403 676
rect 365 524 371 656
rect 317 504 323 516
rect 237 484 243 496
rect 301 464 307 476
rect 45 324 51 356
rect 77 343 83 436
rect 68 337 83 343
rect 61 304 67 316
rect 77 304 83 337
rect 45 284 51 296
rect 93 284 99 376
rect 125 304 131 416
rect 141 304 147 316
rect 221 304 227 436
rect 237 344 243 456
rect 397 424 403 656
rect 125 264 131 296
rect 157 284 163 296
rect 77 124 83 156
rect 109 124 115 236
rect 173 224 179 236
rect 141 144 147 196
rect 205 184 211 276
rect 237 264 243 336
rect 253 284 259 336
rect 269 264 275 356
rect 301 284 307 396
rect 349 344 355 396
rect 381 284 387 316
rect 397 304 403 396
rect 429 263 435 696
rect 445 684 451 716
rect 493 684 499 736
rect 589 724 595 776
rect 525 704 531 716
rect 509 684 515 696
rect 589 684 595 716
rect 621 704 627 836
rect 653 784 659 916
rect 653 704 659 756
rect 621 684 627 696
rect 445 504 451 636
rect 461 564 467 636
rect 525 604 531 676
rect 637 664 643 676
rect 493 504 499 516
rect 509 504 515 556
rect 525 484 531 516
rect 541 504 547 536
rect 605 484 611 576
rect 621 524 627 596
rect 637 564 643 656
rect 653 564 659 636
rect 669 584 675 856
rect 685 844 691 896
rect 781 783 787 936
rect 813 924 819 956
rect 765 777 787 783
rect 685 604 691 716
rect 765 704 771 777
rect 797 743 803 836
rect 829 744 835 836
rect 781 737 803 743
rect 781 724 787 737
rect 781 704 787 716
rect 765 684 771 696
rect 781 684 787 696
rect 829 684 835 696
rect 845 684 851 696
rect 717 584 723 676
rect 733 584 739 636
rect 685 544 691 576
rect 701 544 707 556
rect 765 544 771 576
rect 637 504 643 536
rect 701 524 707 536
rect 717 484 723 496
rect 781 484 787 576
rect 445 304 451 436
rect 461 403 467 436
rect 461 397 483 403
rect 445 264 451 296
rect 413 257 435 263
rect 221 184 227 236
rect 189 104 195 116
rect 221 103 227 176
rect 237 124 243 216
rect 285 164 291 236
rect 349 184 355 236
rect 413 204 419 257
rect 461 243 467 376
rect 477 344 483 397
rect 493 384 499 416
rect 541 344 547 396
rect 477 324 483 336
rect 493 304 499 336
rect 509 304 515 316
rect 541 244 547 336
rect 589 264 595 336
rect 621 304 627 436
rect 685 404 691 476
rect 637 304 643 316
rect 653 304 659 316
rect 621 284 627 296
rect 445 237 467 243
rect 429 224 435 236
rect 445 164 451 237
rect 461 164 467 196
rect 253 124 259 136
rect 285 104 291 116
rect 317 104 323 116
rect 333 104 339 156
rect 365 104 371 136
rect 381 124 387 136
rect 445 124 451 156
rect 525 144 531 176
rect 557 144 563 156
rect 564 137 579 143
rect 509 104 515 116
rect 573 104 579 137
rect 589 124 595 176
rect 653 144 659 256
rect 669 204 675 236
rect 685 164 691 296
rect 701 284 707 396
rect 733 324 739 476
rect 797 384 803 616
rect 829 584 835 596
rect 877 524 883 1037
rect 893 924 899 1016
rect 909 1004 915 1036
rect 941 904 947 956
rect 973 924 979 1016
rect 909 884 915 896
rect 893 724 899 836
rect 925 804 931 836
rect 941 764 947 896
rect 973 783 979 836
rect 973 777 995 783
rect 973 724 979 756
rect 989 704 995 777
rect 893 564 899 696
rect 1005 644 1011 1156
rect 1021 1024 1027 1076
rect 1037 1044 1043 1116
rect 1069 1104 1075 1116
rect 1053 1084 1059 1096
rect 1053 1064 1059 1076
rect 1021 944 1027 996
rect 1037 984 1043 1036
rect 1085 924 1091 1216
rect 1117 1124 1123 1136
rect 1101 904 1107 1036
rect 1149 984 1155 1396
rect 1165 1084 1171 1456
rect 1197 1344 1203 1516
rect 1213 1464 1219 1756
rect 1213 1384 1219 1436
rect 1229 1404 1235 1757
rect 1341 1724 1347 1956
rect 1357 1944 1363 1976
rect 1373 1944 1379 1956
rect 1357 1884 1363 1916
rect 1373 1904 1379 1916
rect 1389 1864 1395 1916
rect 1405 1864 1411 2097
rect 1501 2064 1507 2096
rect 1661 2084 1667 2116
rect 1421 1984 1427 2056
rect 1405 1844 1411 1856
rect 1421 1804 1427 1936
rect 1437 1904 1443 1976
rect 1453 1924 1459 2016
rect 1560 2006 1566 2014
rect 1574 2006 1580 2014
rect 1588 2006 1594 2014
rect 1602 2006 1608 2014
rect 1453 1884 1459 1916
rect 1501 1904 1507 1916
rect 1565 1884 1571 1956
rect 1645 1924 1651 1996
rect 1373 1744 1379 1776
rect 1421 1764 1427 1776
rect 1357 1704 1363 1716
rect 1373 1704 1379 1736
rect 1421 1724 1427 1756
rect 1437 1744 1443 1876
rect 1469 1804 1475 1836
rect 1517 1824 1523 1876
rect 1261 1664 1267 1696
rect 1261 1584 1267 1656
rect 1277 1563 1283 1596
rect 1293 1564 1299 1636
rect 1261 1557 1283 1563
rect 1261 1484 1267 1557
rect 1293 1504 1299 1536
rect 1197 1324 1203 1336
rect 1213 1304 1219 1316
rect 1181 1104 1187 1136
rect 1133 904 1139 916
rect 1149 904 1155 916
rect 1021 784 1027 876
rect 1101 824 1107 896
rect 1165 884 1171 956
rect 1197 944 1203 1236
rect 1261 1184 1267 1476
rect 1277 1444 1283 1476
rect 1293 1324 1299 1376
rect 1213 1004 1219 1036
rect 1197 924 1203 936
rect 1037 684 1043 736
rect 1101 724 1107 796
rect 1133 784 1139 836
rect 1117 724 1123 776
rect 1149 704 1155 796
rect 1165 724 1171 836
rect 1181 704 1187 816
rect 1069 684 1075 696
rect 1213 664 1219 996
rect 1229 924 1235 1136
rect 1261 1104 1267 1176
rect 1309 1124 1315 1496
rect 1325 1463 1331 1656
rect 1341 1504 1347 1576
rect 1357 1504 1363 1656
rect 1389 1644 1395 1716
rect 1325 1457 1347 1463
rect 1325 1324 1331 1436
rect 1341 1344 1347 1457
rect 1357 1404 1363 1476
rect 1389 1363 1395 1636
rect 1405 1484 1411 1636
rect 1453 1564 1459 1796
rect 1533 1744 1539 1836
rect 1469 1684 1475 1696
rect 1501 1663 1507 1736
rect 1485 1657 1507 1663
rect 1517 1717 1532 1723
rect 1485 1504 1491 1657
rect 1501 1584 1507 1636
rect 1517 1624 1523 1717
rect 1549 1704 1555 1776
rect 1549 1684 1555 1696
rect 1533 1604 1539 1636
rect 1560 1606 1566 1614
rect 1574 1606 1580 1614
rect 1588 1606 1594 1614
rect 1602 1606 1608 1614
rect 1549 1504 1555 1516
rect 1405 1424 1411 1456
rect 1421 1404 1427 1436
rect 1437 1424 1443 1476
rect 1380 1357 1395 1363
rect 1469 1324 1475 1376
rect 1533 1324 1539 1476
rect 1565 1324 1571 1556
rect 1581 1364 1587 1456
rect 1597 1344 1603 1476
rect 1629 1384 1635 1796
rect 1661 1744 1667 2016
rect 1677 1983 1683 2036
rect 1693 2024 1699 2476
rect 1725 2384 1731 2436
rect 1837 2384 1843 2436
rect 1709 2284 1715 2336
rect 1725 2304 1731 2356
rect 1773 2284 1779 2356
rect 1853 2344 1859 2356
rect 1805 2264 1811 2336
rect 1837 2304 1843 2336
rect 1725 2204 1731 2236
rect 1869 2224 1875 2496
rect 1917 2484 1923 2556
rect 1997 2544 2003 2596
rect 2013 2564 2019 2636
rect 2045 2584 2051 2856
rect 2077 2704 2083 2836
rect 2109 2784 2115 2896
rect 2141 2883 2147 2896
rect 2173 2884 2179 2916
rect 2237 2897 2252 2903
rect 2125 2877 2147 2883
rect 2125 2724 2131 2877
rect 2141 2784 2147 2856
rect 2173 2764 2179 2836
rect 2237 2744 2243 2897
rect 2301 2864 2307 2916
rect 2285 2744 2291 2756
rect 2132 2717 2147 2723
rect 2141 2664 2147 2717
rect 2189 2704 2195 2736
rect 2205 2704 2211 2716
rect 2221 2704 2227 2736
rect 2173 2684 2179 2696
rect 2237 2664 2243 2736
rect 2317 2724 2323 2936
rect 2349 2904 2355 2936
rect 2381 2884 2387 2956
rect 2381 2764 2387 2836
rect 2285 2684 2291 2696
rect 2301 2684 2307 2696
rect 2317 2664 2323 2716
rect 2333 2704 2339 2756
rect 2413 2744 2419 2836
rect 2445 2824 2451 3056
rect 2509 3024 2515 3036
rect 2477 2964 2483 3016
rect 2557 2984 2563 3176
rect 2589 3104 2595 3236
rect 2605 3184 2611 3276
rect 2685 3264 2691 3316
rect 2717 3264 2723 3296
rect 2605 3104 2611 3156
rect 2637 3144 2643 3156
rect 2685 3144 2691 3236
rect 2733 3184 2739 3457
rect 2749 3324 2755 3356
rect 2765 3344 2771 3396
rect 2813 3324 2819 3356
rect 2829 3344 2835 3396
rect 2861 3384 2867 3436
rect 2893 3384 2899 3436
rect 2781 3284 2787 3296
rect 2589 3084 2595 3096
rect 2669 3084 2675 3116
rect 2573 3004 2579 3036
rect 2493 2904 2499 2956
rect 2541 2924 2547 2936
rect 2525 2884 2531 2916
rect 2589 2904 2595 2976
rect 2621 2924 2627 2996
rect 2685 2984 2691 3116
rect 2701 3104 2707 3176
rect 2749 3164 2755 3236
rect 2813 3144 2819 3276
rect 2653 2944 2659 2956
rect 2701 2924 2707 3096
rect 2717 2904 2723 3116
rect 2813 3084 2819 3136
rect 2845 3124 2851 3316
rect 2877 3144 2883 3336
rect 2861 3104 2867 3136
rect 2877 3104 2883 3136
rect 2749 3064 2755 3076
rect 2733 2944 2739 3036
rect 2797 2964 2803 3036
rect 2813 2984 2819 3036
rect 2772 2917 2812 2923
rect 2573 2897 2588 2903
rect 2429 2724 2435 2756
rect 2445 2664 2451 2716
rect 2461 2704 2467 2736
rect 2573 2704 2579 2897
rect 2477 2684 2483 2696
rect 2500 2657 2508 2663
rect 1981 2504 1987 2536
rect 1997 2524 2003 2536
rect 2013 2524 2019 2536
rect 2077 2504 2083 2556
rect 2109 2544 2115 2576
rect 2125 2524 2131 2556
rect 1901 2364 1907 2436
rect 1949 2404 1955 2436
rect 1965 2344 1971 2456
rect 1997 2384 2003 2476
rect 1885 2304 1891 2316
rect 1709 2084 1715 2116
rect 1725 2064 1731 2116
rect 1757 2104 1763 2156
rect 1901 2144 1907 2296
rect 1933 2264 1939 2316
rect 1981 2304 1987 2356
rect 1997 2324 2003 2376
rect 2061 2324 2067 2396
rect 2045 2284 2051 2316
rect 2093 2284 2099 2376
rect 2141 2344 2147 2656
rect 2157 2504 2163 2536
rect 2173 2483 2179 2656
rect 2205 2484 2211 2516
rect 2237 2504 2243 2616
rect 2269 2524 2275 2636
rect 2365 2584 2371 2636
rect 2301 2544 2307 2576
rect 2317 2524 2323 2556
rect 2157 2477 2179 2483
rect 2157 2304 2163 2477
rect 2189 2464 2195 2476
rect 2173 2404 2179 2436
rect 2205 2364 2211 2476
rect 2253 2444 2259 2516
rect 2269 2484 2275 2516
rect 2333 2464 2339 2516
rect 2365 2503 2371 2556
rect 2397 2504 2403 2616
rect 2413 2524 2419 2536
rect 2356 2497 2371 2503
rect 2349 2444 2355 2496
rect 2429 2484 2435 2516
rect 2461 2484 2467 2556
rect 2493 2504 2499 2656
rect 2525 2644 2531 2676
rect 2621 2664 2627 2716
rect 2589 2644 2595 2656
rect 2525 2544 2531 2636
rect 2621 2624 2627 2656
rect 2637 2584 2643 2816
rect 2653 2644 2659 2776
rect 2701 2724 2707 2896
rect 2749 2884 2755 2916
rect 2717 2724 2723 2816
rect 2749 2784 2755 2856
rect 2669 2704 2675 2716
rect 2685 2664 2691 2676
rect 2653 2524 2659 2536
rect 2669 2504 2675 2536
rect 2269 2384 2275 2416
rect 2116 2257 2131 2263
rect 1949 2184 1955 2236
rect 1965 2144 1971 2156
rect 1997 2144 2003 2196
rect 2029 2164 2035 2236
rect 1805 2084 1811 2116
rect 1821 2084 1827 2136
rect 1869 2084 1875 2116
rect 1885 2084 1891 2136
rect 1917 2084 1923 2136
rect 1997 2104 2003 2136
rect 2013 2124 2019 2156
rect 2061 2144 2067 2236
rect 2125 2144 2131 2257
rect 2173 2184 2179 2276
rect 2061 2084 2067 2136
rect 2125 2124 2131 2136
rect 2141 2124 2147 2176
rect 2173 2124 2179 2176
rect 2189 2164 2195 2296
rect 2237 2244 2243 2316
rect 2349 2304 2355 2396
rect 2365 2344 2371 2436
rect 2269 2284 2275 2296
rect 2365 2284 2371 2316
rect 2413 2304 2419 2316
rect 2253 2244 2259 2256
rect 2301 2164 2307 2236
rect 2317 2204 2323 2276
rect 2429 2264 2435 2316
rect 2477 2304 2483 2316
rect 2157 2104 2163 2116
rect 2189 2084 2195 2156
rect 2253 2104 2259 2116
rect 2269 2104 2275 2116
rect 2253 2084 2259 2096
rect 2237 2064 2243 2076
rect 2301 2064 2307 2116
rect 1677 1977 1699 1983
rect 1677 1884 1683 1956
rect 1693 1884 1699 1977
rect 1725 1964 1731 2036
rect 1741 1904 1747 1916
rect 1757 1884 1763 1896
rect 1773 1824 1779 1936
rect 1805 1924 1811 2036
rect 1869 2004 1875 2036
rect 1901 1924 1907 2056
rect 1805 1884 1811 1896
rect 1821 1824 1827 1876
rect 1869 1864 1875 1896
rect 1949 1884 1955 1996
rect 1965 1904 1971 2036
rect 2013 1924 2019 2036
rect 2093 2004 2099 2036
rect 2045 1944 2051 1956
rect 2061 1944 2067 1956
rect 2077 1924 2083 1976
rect 2093 1904 2099 1956
rect 2109 1884 2115 1896
rect 2141 1864 2147 1976
rect 2221 1964 2227 2036
rect 2205 1884 2211 1916
rect 2221 1904 2227 1936
rect 2237 1904 2243 2016
rect 2317 1904 2323 2196
rect 2413 2184 2419 2216
rect 2365 2124 2371 2136
rect 2349 2084 2355 2116
rect 2333 2024 2339 2036
rect 2381 1984 2387 2076
rect 2397 2044 2403 2156
rect 2413 2024 2419 2096
rect 2429 2064 2435 2256
rect 2493 2224 2499 2496
rect 2557 2484 2563 2496
rect 2525 2464 2531 2476
rect 2573 2464 2579 2476
rect 2509 2304 2515 2436
rect 2573 2424 2579 2436
rect 2589 2384 2595 2476
rect 2605 2343 2611 2456
rect 2653 2443 2659 2496
rect 2685 2483 2691 2636
rect 2701 2604 2707 2696
rect 2701 2524 2707 2576
rect 2733 2544 2739 2756
rect 2749 2704 2755 2756
rect 2749 2584 2755 2676
rect 2628 2437 2659 2443
rect 2669 2477 2691 2483
rect 2669 2384 2675 2477
rect 2717 2384 2723 2456
rect 2605 2337 2627 2343
rect 2605 2264 2611 2316
rect 2621 2304 2627 2337
rect 2685 2304 2691 2336
rect 2701 2304 2707 2376
rect 2749 2363 2755 2576
rect 2765 2384 2771 2876
rect 2797 2844 2803 2876
rect 2845 2784 2851 3056
rect 2877 2984 2883 3076
rect 2861 2944 2867 2976
rect 2893 2964 2899 3136
rect 2909 3124 2915 3156
rect 2909 3044 2915 3116
rect 2925 3004 2931 3216
rect 2941 3184 2947 3436
rect 2957 3404 2963 3436
rect 2973 3284 2979 3316
rect 2989 3304 2995 3436
rect 2957 3264 2963 3276
rect 2941 3064 2947 3096
rect 2909 2944 2915 2976
rect 2861 2744 2867 2776
rect 2877 2724 2883 2896
rect 2893 2864 2899 2936
rect 2925 2923 2931 2976
rect 2957 2963 2963 3116
rect 2916 2917 2931 2923
rect 2941 2957 2963 2963
rect 2909 2904 2915 2916
rect 2900 2857 2915 2863
rect 2909 2763 2915 2857
rect 2925 2784 2931 2816
rect 2909 2757 2931 2763
rect 2813 2703 2819 2716
rect 2813 2697 2828 2703
rect 2829 2684 2835 2696
rect 2845 2684 2851 2696
rect 2788 2677 2796 2683
rect 2781 2584 2787 2656
rect 2781 2564 2787 2576
rect 2797 2544 2803 2556
rect 2829 2504 2835 2636
rect 2845 2544 2851 2676
rect 2861 2484 2867 2636
rect 2749 2357 2771 2363
rect 2724 2337 2748 2343
rect 2765 2323 2771 2357
rect 2749 2317 2771 2323
rect 2477 2104 2483 2156
rect 2509 2144 2515 2196
rect 2573 2164 2579 2176
rect 2445 1984 2451 2016
rect 2493 1984 2499 2036
rect 2525 1984 2531 2136
rect 2557 2084 2563 2096
rect 2237 1884 2243 1896
rect 2333 1884 2339 1936
rect 2365 1883 2371 1936
rect 2397 1924 2403 1936
rect 2461 1904 2467 1916
rect 2388 1897 2444 1903
rect 2365 1877 2387 1883
rect 2269 1864 2275 1876
rect 2276 1857 2291 1863
rect 2285 1844 2291 1857
rect 1709 1744 1715 1756
rect 1725 1744 1731 1776
rect 1997 1764 2003 1776
rect 1773 1744 1779 1756
rect 1652 1717 1667 1723
rect 1645 1464 1651 1656
rect 1661 1584 1667 1717
rect 1693 1683 1699 1736
rect 1709 1704 1715 1736
rect 1885 1724 1891 1736
rect 1853 1717 1868 1723
rect 1789 1684 1795 1716
rect 1693 1677 1715 1683
rect 1661 1524 1667 1576
rect 1709 1484 1715 1677
rect 1837 1664 1843 1696
rect 1853 1644 1859 1717
rect 1933 1704 1939 1716
rect 1789 1523 1795 1636
rect 1780 1517 1795 1523
rect 1725 1484 1731 1496
rect 1661 1444 1667 1476
rect 1709 1464 1715 1476
rect 1389 1264 1395 1296
rect 1533 1284 1539 1296
rect 1549 1284 1555 1316
rect 1565 1304 1571 1316
rect 1261 1044 1267 1076
rect 1229 904 1235 916
rect 1293 863 1299 1076
rect 1309 1004 1315 1096
rect 1325 983 1331 1196
rect 1341 1064 1347 1236
rect 1389 1224 1395 1256
rect 1597 1244 1603 1336
rect 1677 1304 1683 1376
rect 1709 1364 1715 1456
rect 1741 1364 1747 1376
rect 1693 1344 1699 1356
rect 1773 1344 1779 1356
rect 1821 1344 1827 1596
rect 1853 1504 1859 1556
rect 1901 1504 1907 1636
rect 1917 1564 1923 1676
rect 1933 1524 1939 1536
rect 1837 1484 1843 1496
rect 1901 1464 1907 1476
rect 1917 1384 1923 1496
rect 1965 1484 1971 1716
rect 2013 1704 2019 1756
rect 2045 1724 2051 1836
rect 2061 1744 2067 1776
rect 2125 1764 2131 1836
rect 2125 1704 2131 1736
rect 2157 1704 2163 1736
rect 2173 1724 2179 1836
rect 2237 1724 2243 1756
rect 2253 1744 2259 1836
rect 2045 1624 2051 1636
rect 1997 1484 2003 1536
rect 2013 1464 2019 1480
rect 1885 1357 1932 1363
rect 1613 1264 1619 1296
rect 1773 1284 1779 1336
rect 1805 1304 1811 1316
rect 1853 1303 1859 1356
rect 1885 1344 1891 1357
rect 1949 1344 1955 1456
rect 1965 1384 1971 1436
rect 1997 1364 2003 1376
rect 2013 1344 2019 1356
rect 1844 1297 1859 1303
rect 1837 1264 1843 1296
rect 1629 1244 1635 1256
rect 1357 1064 1363 1116
rect 1405 1104 1411 1156
rect 1421 1104 1427 1236
rect 1437 1144 1443 1156
rect 1469 1144 1475 1236
rect 1517 1164 1523 1236
rect 1560 1206 1566 1214
rect 1574 1206 1580 1214
rect 1588 1206 1594 1214
rect 1602 1206 1608 1214
rect 1565 1124 1571 1176
rect 1597 1104 1603 1136
rect 1421 1083 1427 1096
rect 1613 1084 1619 1096
rect 1412 1077 1427 1083
rect 1629 1083 1635 1236
rect 1741 1184 1747 1196
rect 1757 1184 1763 1236
rect 1869 1184 1875 1256
rect 1620 1077 1635 1083
rect 1645 1064 1651 1176
rect 1821 1144 1827 1156
rect 1757 1117 1772 1123
rect 1709 1064 1715 1116
rect 1725 1104 1731 1116
rect 1309 977 1331 983
rect 1309 964 1315 977
rect 1309 944 1315 956
rect 1277 857 1299 863
rect 1229 724 1235 776
rect 1229 704 1235 716
rect 1261 704 1267 716
rect 1277 684 1283 857
rect 1325 844 1331 956
rect 1341 904 1347 1056
rect 1357 944 1363 1056
rect 1517 1024 1523 1036
rect 1405 904 1411 976
rect 1501 964 1507 976
rect 1421 904 1427 916
rect 1389 864 1395 876
rect 1293 744 1299 836
rect 1421 784 1427 896
rect 1437 884 1443 916
rect 1453 864 1459 876
rect 1565 844 1571 936
rect 1613 864 1619 916
rect 1629 884 1635 936
rect 1293 664 1299 676
rect 893 524 899 536
rect 813 497 828 503
rect 765 324 771 356
rect 637 124 643 136
rect 653 124 659 136
rect 212 97 227 103
rect 605 84 611 96
rect 717 84 723 296
rect 781 284 787 356
rect 813 344 819 497
rect 861 464 867 516
rect 909 444 915 636
rect 925 524 931 636
rect 957 524 963 636
rect 957 504 963 516
rect 829 324 835 416
rect 925 404 931 436
rect 845 384 851 396
rect 909 304 915 316
rect 749 264 755 276
rect 797 244 803 296
rect 861 264 867 276
rect 909 224 915 276
rect 925 244 931 396
rect 973 323 979 556
rect 1005 524 1011 596
rect 1069 524 1075 596
rect 1117 584 1123 636
rect 1213 584 1219 636
rect 1229 564 1235 636
rect 1309 624 1315 756
rect 1373 704 1379 736
rect 1341 664 1347 676
rect 1389 664 1395 676
rect 1325 584 1331 636
rect 1357 584 1363 616
rect 989 464 995 476
rect 1005 464 1011 476
rect 989 344 995 456
rect 1021 384 1027 496
rect 1053 464 1059 476
rect 1021 324 1027 336
rect 1037 324 1043 396
rect 1069 344 1075 436
rect 1085 364 1091 496
rect 1117 424 1123 516
rect 1133 484 1139 536
rect 1165 524 1171 556
rect 1245 503 1251 516
rect 1245 497 1260 503
rect 1133 384 1139 396
rect 1245 384 1251 497
rect 1277 424 1283 516
rect 1293 484 1299 536
rect 1325 384 1331 516
rect 1341 484 1347 556
rect 1405 543 1411 636
rect 1421 584 1427 716
rect 1437 563 1443 836
rect 1517 784 1523 836
rect 1560 806 1566 814
rect 1574 806 1580 814
rect 1588 806 1594 814
rect 1602 806 1608 814
rect 1661 784 1667 856
rect 1469 704 1475 736
rect 1453 684 1459 696
rect 1453 664 1459 676
rect 1533 663 1539 716
rect 1693 664 1699 836
rect 1709 684 1715 976
rect 1725 944 1731 1056
rect 1725 904 1731 916
rect 1741 884 1747 936
rect 1757 764 1763 1117
rect 1773 1104 1779 1116
rect 1805 1044 1811 1136
rect 1821 1124 1827 1136
rect 1821 1024 1827 1096
rect 1837 964 1843 1156
rect 1901 1144 1907 1336
rect 2029 1324 2035 1576
rect 2061 1504 2067 1516
rect 2093 1504 2099 1676
rect 2109 1664 2115 1696
rect 2125 1684 2131 1696
rect 2141 1464 2147 1476
rect 2157 1464 2163 1656
rect 2189 1604 2195 1696
rect 2045 1323 2051 1436
rect 2125 1404 2131 1436
rect 2109 1364 2115 1376
rect 2173 1364 2179 1516
rect 2205 1504 2211 1696
rect 2269 1584 2275 1836
rect 2301 1683 2307 1876
rect 2301 1677 2323 1683
rect 2317 1584 2323 1677
rect 2333 1584 2339 1856
rect 2365 1784 2371 1816
rect 2381 1804 2387 1877
rect 2365 1724 2371 1736
rect 2365 1684 2371 1716
rect 2381 1644 2387 1696
rect 2397 1644 2403 1897
rect 2477 1804 2483 1936
rect 2541 1904 2547 1936
rect 2493 1824 2499 1896
rect 2541 1803 2547 1896
rect 2557 1824 2563 1876
rect 2573 1804 2579 2076
rect 2589 1984 2595 2116
rect 2605 2064 2611 2136
rect 2621 2097 2636 2103
rect 2621 1984 2627 2097
rect 2637 2084 2643 2096
rect 2653 1943 2659 2236
rect 2669 2184 2675 2256
rect 2717 2244 2723 2316
rect 2749 2184 2755 2317
rect 2781 2264 2787 2456
rect 2829 2383 2835 2476
rect 2845 2404 2851 2436
rect 2893 2404 2899 2756
rect 2909 2724 2915 2736
rect 2925 2704 2931 2757
rect 2941 2724 2947 2957
rect 2957 2743 2963 2816
rect 2973 2763 2979 2996
rect 2989 2964 2995 3296
rect 3005 3284 3011 3336
rect 3021 3304 3027 3436
rect 3037 3384 3043 3517
rect 3037 3264 3043 3296
rect 3037 3184 3043 3256
rect 3069 3164 3075 3516
rect 3085 3464 3091 3496
rect 3117 3484 3123 3636
rect 3197 3544 3203 3636
rect 3229 3584 3235 3616
rect 3213 3504 3219 3516
rect 3213 3484 3219 3496
rect 3245 3424 3251 3516
rect 3261 3504 3267 3736
rect 3277 3704 3283 3716
rect 3293 3704 3299 3736
rect 3277 3524 3283 3696
rect 3325 3584 3331 3757
rect 3341 3704 3347 3736
rect 3357 3604 3363 3736
rect 3389 3704 3395 3936
rect 3501 3924 3507 4157
rect 3517 4124 3523 4156
rect 3549 4144 3555 4156
rect 3565 4144 3571 4176
rect 3581 4123 3587 4197
rect 3597 4184 3603 4456
rect 3645 4384 3651 4536
rect 3613 4184 3619 4276
rect 3629 4144 3635 4236
rect 3645 4224 3651 4256
rect 3645 4144 3651 4216
rect 3572 4117 3587 4123
rect 3437 3904 3443 3916
rect 3405 3644 3411 3896
rect 3421 3824 3427 3896
rect 3437 3764 3443 3836
rect 3453 3784 3459 3816
rect 3501 3744 3507 3916
rect 3517 3904 3523 3916
rect 3517 3784 3523 3896
rect 3533 3744 3539 4016
rect 3581 3904 3587 3976
rect 3549 3784 3555 3896
rect 3597 3884 3603 3936
rect 3581 3784 3587 3856
rect 3597 3764 3603 3836
rect 3613 3824 3619 4136
rect 3661 4124 3667 4296
rect 3693 4184 3699 4336
rect 3709 4244 3715 4316
rect 3725 4304 3731 4516
rect 3741 4464 3747 4536
rect 3805 4384 3811 4496
rect 3869 4384 3875 4396
rect 3741 4184 3747 4296
rect 3789 4284 3795 4336
rect 3805 4184 3811 4276
rect 3821 4264 3827 4316
rect 3837 4184 3843 4296
rect 3901 4244 3907 4516
rect 3933 4504 3939 4536
rect 3917 4324 3923 4436
rect 3933 4404 3939 4496
rect 3949 4384 3955 4476
rect 3997 4444 4003 4516
rect 4029 4323 4035 4536
rect 4061 4384 4067 4576
rect 4157 4564 4163 4896
rect 4397 4884 4403 4916
rect 4429 4904 4435 4956
rect 4445 4904 4451 4956
rect 4413 4864 4419 4876
rect 4301 4744 4307 4756
rect 4365 4744 4371 4756
rect 4237 4684 4243 4736
rect 4173 4584 4179 4676
rect 4237 4584 4243 4676
rect 4253 4644 4259 4696
rect 4269 4664 4275 4716
rect 4317 4704 4323 4736
rect 4333 4704 4339 4716
rect 4381 4704 4387 4736
rect 4397 4724 4403 4736
rect 4413 4704 4419 4716
rect 4285 4584 4291 4596
rect 4381 4584 4387 4676
rect 4429 4664 4435 4896
rect 4141 4504 4147 4516
rect 4077 4444 4083 4496
rect 4125 4384 4131 4456
rect 4020 4317 4035 4323
rect 3709 4104 3715 4136
rect 3741 4104 3747 4136
rect 3677 3944 3683 3976
rect 3645 3863 3651 3916
rect 3661 3904 3667 3936
rect 3709 3903 3715 4096
rect 3741 3984 3747 4076
rect 3757 4044 3763 4136
rect 3773 4124 3779 4156
rect 3789 3964 3795 4116
rect 3853 4104 3859 4236
rect 3917 4184 3923 4316
rect 3965 4284 3971 4316
rect 3805 4084 3811 4096
rect 3725 3924 3731 3936
rect 3741 3904 3747 3956
rect 3709 3897 3731 3903
rect 3636 3857 3651 3863
rect 3645 3784 3651 3857
rect 3693 3784 3699 3816
rect 3709 3764 3715 3836
rect 3725 3784 3731 3897
rect 3757 3824 3763 3916
rect 3773 3904 3779 3916
rect 3789 3884 3795 3956
rect 3613 3744 3619 3756
rect 3453 3737 3468 3743
rect 3357 3584 3363 3596
rect 3112 3406 3118 3414
rect 3126 3406 3132 3414
rect 3140 3406 3146 3414
rect 3154 3406 3160 3414
rect 3213 3384 3219 3416
rect 3197 3364 3203 3376
rect 3229 3344 3235 3356
rect 3149 3324 3155 3336
rect 3229 3324 3235 3336
rect 3181 3283 3187 3316
rect 3245 3303 3251 3416
rect 3261 3344 3267 3416
rect 3277 3384 3283 3436
rect 3309 3384 3315 3536
rect 3325 3424 3331 3496
rect 3341 3464 3347 3476
rect 3245 3297 3260 3303
rect 3165 3277 3187 3283
rect 3165 3184 3171 3277
rect 3213 3184 3219 3276
rect 3293 3264 3299 3336
rect 3309 3184 3315 3316
rect 3325 3304 3331 3356
rect 3341 3344 3347 3416
rect 3357 3364 3363 3516
rect 3389 3484 3395 3496
rect 3373 3344 3379 3356
rect 3005 3104 3011 3116
rect 3021 3084 3027 3116
rect 3037 3104 3043 3116
rect 3005 2964 3011 3016
rect 3005 2924 3011 2936
rect 2989 2904 2995 2916
rect 2989 2884 2995 2896
rect 3021 2884 3027 3076
rect 3037 3004 3043 3096
rect 3053 2924 3059 3136
rect 3069 2944 3075 3156
rect 3085 2944 3091 3096
rect 3165 3044 3171 3076
rect 3112 3006 3118 3014
rect 3126 3006 3132 3014
rect 3140 3006 3146 3014
rect 3154 3006 3160 3014
rect 3181 3004 3187 3136
rect 3197 3084 3203 3156
rect 3213 3064 3219 3096
rect 3213 2984 3219 3056
rect 3204 2957 3219 2963
rect 3213 2944 3219 2957
rect 2989 2784 2995 2816
rect 2973 2757 2995 2763
rect 2957 2737 2972 2743
rect 2989 2724 2995 2757
rect 2941 2644 2947 2716
rect 2989 2644 2995 2696
rect 2941 2504 2947 2596
rect 2973 2524 2979 2616
rect 3037 2584 3043 2896
rect 3053 2864 3059 2916
rect 3069 2884 3075 2916
rect 3085 2904 3091 2936
rect 3149 2904 3155 2936
rect 3181 2904 3187 2936
rect 3213 2904 3219 2916
rect 3053 2664 3059 2716
rect 3069 2644 3075 2856
rect 3085 2844 3091 2896
rect 3181 2837 3219 2843
rect 3085 2744 3091 2816
rect 3101 2784 3107 2836
rect 2989 2524 2995 2556
rect 2909 2484 2915 2496
rect 2989 2484 2995 2516
rect 3021 2504 3027 2556
rect 2829 2377 2899 2383
rect 2797 2337 2812 2343
rect 2797 2324 2803 2337
rect 2829 2323 2835 2377
rect 2845 2357 2883 2363
rect 2845 2344 2851 2357
rect 2861 2323 2867 2336
rect 2829 2317 2867 2323
rect 2813 2264 2819 2316
rect 2877 2304 2883 2357
rect 2893 2344 2899 2377
rect 2845 2284 2851 2296
rect 2813 2244 2819 2256
rect 2685 2024 2691 2136
rect 2733 2084 2739 2096
rect 2797 2064 2803 2136
rect 2644 1937 2659 1943
rect 2605 1863 2611 1916
rect 2701 1904 2707 2036
rect 2717 2024 2723 2036
rect 2717 1944 2723 2016
rect 2813 1964 2819 2076
rect 2765 1944 2771 1956
rect 2733 1924 2739 1936
rect 2596 1857 2611 1863
rect 2621 1824 2627 1896
rect 2685 1884 2691 1896
rect 2701 1884 2707 1896
rect 2541 1797 2563 1803
rect 2445 1784 2451 1796
rect 2557 1784 2563 1797
rect 2477 1724 2483 1776
rect 2413 1684 2419 1716
rect 2445 1683 2451 1716
rect 2525 1704 2531 1756
rect 2589 1724 2595 1736
rect 2605 1704 2611 1716
rect 2445 1677 2460 1683
rect 2621 1664 2627 1736
rect 2637 1724 2643 1796
rect 2717 1764 2723 1916
rect 2733 1844 2739 1916
rect 2381 1584 2387 1596
rect 2637 1584 2643 1656
rect 2669 1624 2675 1696
rect 2701 1684 2707 1736
rect 2717 1704 2723 1716
rect 2733 1704 2739 1756
rect 2749 1704 2755 1716
rect 2189 1464 2195 1496
rect 2205 1444 2211 1456
rect 2221 1384 2227 1576
rect 2237 1444 2243 1456
rect 2253 1404 2259 1456
rect 2269 1384 2275 1436
rect 2045 1317 2060 1323
rect 1933 1144 1939 1196
rect 1949 1184 1955 1316
rect 1965 1163 1971 1276
rect 1956 1157 1971 1163
rect 1853 1024 1859 1116
rect 1949 1104 1955 1136
rect 1885 984 1891 1096
rect 1965 1084 1971 1116
rect 1805 884 1811 916
rect 1821 884 1827 956
rect 1773 704 1779 836
rect 1524 657 1539 663
rect 1597 584 1603 616
rect 1741 584 1747 676
rect 1437 557 1452 563
rect 1389 537 1411 543
rect 1357 524 1363 536
rect 1357 484 1363 516
rect 1341 464 1347 476
rect 1373 464 1379 496
rect 1389 444 1395 537
rect 1405 444 1411 516
rect 1421 484 1427 556
rect 1373 344 1379 356
rect 964 317 979 323
rect 957 304 963 316
rect 989 304 995 316
rect 973 224 979 276
rect 1005 243 1011 316
rect 1053 264 1059 296
rect 989 237 1011 243
rect 861 184 867 196
rect 989 164 995 237
rect 1005 184 1011 216
rect 733 124 739 136
rect 797 124 803 156
rect 813 144 819 156
rect 749 104 755 116
rect 733 64 739 96
rect 877 84 883 96
rect 909 84 915 116
rect 957 84 963 156
rect 1005 143 1011 156
rect 1021 144 1027 236
rect 1101 164 1107 276
rect 1117 184 1123 256
rect 1149 224 1155 316
rect 1229 224 1235 316
rect 1245 284 1251 296
rect 1261 244 1267 336
rect 1325 323 1331 336
rect 1309 317 1331 323
rect 1309 284 1315 317
rect 1389 304 1395 336
rect 1421 324 1427 456
rect 1437 344 1443 536
rect 1485 524 1491 536
rect 1469 463 1475 516
rect 1469 457 1491 463
rect 1469 384 1475 436
rect 1485 364 1491 457
rect 1501 404 1507 516
rect 1533 384 1539 556
rect 1613 524 1619 576
rect 1549 504 1555 516
rect 1629 464 1635 556
rect 1773 544 1779 636
rect 1805 584 1811 796
rect 1837 784 1843 896
rect 1869 844 1875 876
rect 1885 823 1891 896
rect 1869 817 1891 823
rect 1869 764 1875 817
rect 1901 784 1907 1056
rect 1949 984 1955 1036
rect 1981 984 1987 1316
rect 1997 1124 2003 1136
rect 2013 1124 2019 1256
rect 2045 1243 2051 1296
rect 2029 1237 2051 1243
rect 2029 1144 2035 1237
rect 2141 1224 2147 1296
rect 2077 1184 2083 1216
rect 2141 1144 2147 1156
rect 2013 1084 2019 1096
rect 1949 904 1955 916
rect 1965 904 1971 956
rect 1821 724 1827 736
rect 1837 684 1843 696
rect 1869 584 1875 756
rect 1885 744 1891 776
rect 1901 684 1907 696
rect 1917 604 1923 716
rect 1933 584 1939 876
rect 1949 844 1955 876
rect 1965 844 1971 896
rect 1949 784 1955 836
rect 1981 784 1987 916
rect 1997 904 2003 936
rect 2013 804 2019 1076
rect 2061 1004 2067 1136
rect 2077 1104 2083 1136
rect 2157 1124 2163 1296
rect 2173 1184 2179 1296
rect 2189 1204 2195 1316
rect 2205 1244 2211 1336
rect 2237 1304 2243 1356
rect 2253 1324 2259 1336
rect 2189 1144 2195 1196
rect 2141 1104 2147 1116
rect 2045 864 2051 936
rect 2061 843 2067 996
rect 2141 984 2147 1076
rect 2093 904 2099 936
rect 2109 864 2115 916
rect 2116 857 2131 863
rect 2045 837 2067 843
rect 2029 784 2035 796
rect 1949 644 1955 696
rect 1965 584 1971 736
rect 1741 504 1747 516
rect 1757 464 1763 496
rect 1773 484 1779 516
rect 1789 504 1795 536
rect 1821 464 1827 556
rect 1560 406 1566 414
rect 1574 406 1580 414
rect 1588 406 1594 414
rect 1602 406 1608 414
rect 1645 384 1651 396
rect 1373 284 1379 296
rect 996 137 1011 143
rect 1101 104 1107 156
rect 1149 124 1155 156
rect 1165 144 1171 176
rect 1261 144 1267 216
rect 1277 184 1283 236
rect 1325 184 1331 276
rect 1373 164 1379 276
rect 1389 184 1395 236
rect 1421 204 1427 316
rect 1453 264 1459 336
rect 1485 304 1491 316
rect 1501 224 1507 296
rect 1485 184 1491 196
rect 1309 144 1315 156
rect 1405 144 1411 156
rect 1229 104 1235 136
rect 1117 84 1123 96
rect 845 64 851 76
rect 925 64 931 76
rect 1213 -23 1219 -17
rect 1261 -23 1267 -17
rect 1309 -23 1315 -17
rect 1341 -23 1347 136
rect 1357 104 1363 116
rect 1357 -17 1363 96
rect 1357 -23 1379 -17
rect 1437 -23 1443 136
rect 1517 124 1523 336
rect 1565 204 1571 296
rect 1597 224 1603 316
rect 1613 304 1619 356
rect 1677 344 1683 356
rect 1709 324 1715 456
rect 1789 304 1795 316
rect 1693 264 1699 296
rect 1725 264 1731 276
rect 1565 164 1571 196
rect 1725 144 1731 236
rect 1789 224 1795 256
rect 1741 144 1747 196
rect 1805 184 1811 416
rect 1837 404 1843 516
rect 1853 444 1859 536
rect 1885 484 1891 556
rect 1981 523 1987 696
rect 1997 544 2003 616
rect 2013 584 2019 736
rect 2029 644 2035 696
rect 2013 524 2019 576
rect 2029 544 2035 636
rect 2045 584 2051 837
rect 2109 784 2115 836
rect 2061 564 2067 716
rect 2077 564 2083 696
rect 2109 584 2115 676
rect 2125 664 2131 857
rect 2157 784 2163 1116
rect 2205 1104 2211 1236
rect 2221 1144 2227 1196
rect 2237 1144 2243 1276
rect 2269 1244 2275 1316
rect 2285 1184 2291 1536
rect 2301 1504 2307 1536
rect 2365 1504 2371 1536
rect 2397 1524 2403 1556
rect 2701 1544 2707 1676
rect 2717 1624 2723 1636
rect 2733 1564 2739 1696
rect 2381 1504 2387 1516
rect 2317 1484 2323 1496
rect 2365 1384 2371 1496
rect 2397 1443 2403 1516
rect 2413 1484 2419 1516
rect 2429 1504 2435 1516
rect 2541 1504 2547 1516
rect 2589 1504 2595 1516
rect 2381 1437 2403 1443
rect 2317 1304 2323 1376
rect 2253 1124 2259 1136
rect 2173 1044 2179 1076
rect 2237 1004 2243 1116
rect 2253 1104 2259 1116
rect 2301 1084 2307 1236
rect 2317 1144 2323 1276
rect 2333 1184 2339 1376
rect 2349 1184 2355 1236
rect 2381 1184 2387 1437
rect 2397 1344 2403 1356
rect 2397 1224 2403 1316
rect 2413 1284 2419 1436
rect 2429 1384 2435 1496
rect 2621 1484 2627 1536
rect 2644 1497 2652 1503
rect 2717 1503 2723 1536
rect 2765 1523 2771 1896
rect 2813 1824 2819 1836
rect 2765 1517 2787 1523
rect 2708 1497 2723 1503
rect 2477 1444 2483 1456
rect 2509 1444 2515 1476
rect 2477 1364 2483 1396
rect 2493 1384 2499 1416
rect 2525 1364 2531 1436
rect 2557 1424 2563 1476
rect 2429 1204 2435 1276
rect 2349 1124 2355 1136
rect 2333 1104 2339 1116
rect 2349 1064 2355 1116
rect 2365 1043 2371 1116
rect 2381 1084 2387 1096
rect 2381 1044 2387 1076
rect 2349 1037 2371 1043
rect 2269 924 2275 1016
rect 2189 884 2195 916
rect 2221 904 2227 916
rect 2333 884 2339 896
rect 2173 844 2179 876
rect 2189 784 2195 816
rect 2157 664 2163 696
rect 2173 684 2179 696
rect 2125 637 2140 643
rect 2125 564 2131 637
rect 2141 564 2147 616
rect 2157 584 2163 656
rect 2093 544 2099 556
rect 1965 517 1987 523
rect 1965 504 1971 517
rect 1901 444 1907 496
rect 1933 384 1939 456
rect 2029 384 2035 476
rect 2077 384 2083 516
rect 2157 504 2163 576
rect 2189 524 2195 696
rect 2205 664 2211 756
rect 2253 744 2259 836
rect 2349 764 2355 1037
rect 2397 1003 2403 1156
rect 2445 1144 2451 1296
rect 2477 1184 2483 1316
rect 2525 1264 2531 1316
rect 2541 1304 2547 1396
rect 2557 1324 2563 1336
rect 2573 1264 2579 1276
rect 2381 997 2403 1003
rect 2381 924 2387 997
rect 2413 924 2419 976
rect 2429 944 2435 1076
rect 2445 1044 2451 1096
rect 2461 924 2467 936
rect 2381 863 2387 916
rect 2493 884 2499 1196
rect 2509 1104 2515 1216
rect 2605 1184 2611 1336
rect 2621 1304 2627 1316
rect 2621 1164 2627 1256
rect 2637 1183 2643 1436
rect 2653 1384 2659 1476
rect 2717 1464 2723 1476
rect 2692 1457 2707 1463
rect 2685 1384 2691 1436
rect 2701 1384 2707 1457
rect 2701 1224 2707 1336
rect 2637 1177 2659 1183
rect 2509 1084 2515 1096
rect 2525 1024 2531 1036
rect 2557 1004 2563 1056
rect 2509 924 2515 956
rect 2541 924 2547 976
rect 2365 857 2387 863
rect 2365 824 2371 857
rect 2381 784 2387 836
rect 2429 764 2435 836
rect 2269 544 2275 676
rect 2317 624 2323 716
rect 2461 704 2467 776
rect 2493 744 2499 836
rect 2493 723 2499 736
rect 2525 724 2531 896
rect 2541 884 2547 896
rect 2573 883 2579 1076
rect 2589 1064 2595 1116
rect 2637 1104 2643 1156
rect 2653 1144 2659 1177
rect 2669 1104 2675 1156
rect 2685 1104 2691 1116
rect 2733 1104 2739 1436
rect 2749 1264 2755 1476
rect 2765 1384 2771 1456
rect 2765 1304 2771 1316
rect 2781 1304 2787 1517
rect 2797 1464 2803 1696
rect 2813 1684 2819 1696
rect 2829 1663 2835 2256
rect 2845 2084 2851 2136
rect 2845 2064 2851 2076
rect 2845 1924 2851 1936
rect 2861 1884 2867 2296
rect 2909 2284 2915 2296
rect 2925 2204 2931 2396
rect 2941 2384 2947 2476
rect 2957 2437 2972 2443
rect 2957 2324 2963 2437
rect 2973 2384 2979 2416
rect 3005 2324 3011 2416
rect 2877 1904 2883 2176
rect 2941 2144 2947 2296
rect 2957 2184 2963 2276
rect 2973 2244 2979 2316
rect 3021 2304 3027 2476
rect 3069 2444 3075 2516
rect 3085 2444 3091 2716
rect 3117 2703 3123 2816
rect 3181 2784 3187 2837
rect 3213 2824 3219 2837
rect 3197 2784 3203 2816
rect 3165 2724 3171 2756
rect 3181 2724 3187 2756
rect 3213 2724 3219 2776
rect 3229 2764 3235 3136
rect 3245 3104 3251 3116
rect 3245 2984 3251 3096
rect 3277 3064 3283 3116
rect 3245 2783 3251 2956
rect 3261 2904 3267 2996
rect 3277 2864 3283 2996
rect 3293 2944 3299 3136
rect 3357 3064 3363 3336
rect 3373 3304 3379 3336
rect 3405 3323 3411 3536
rect 3421 3364 3427 3736
rect 3437 3584 3443 3636
rect 3453 3524 3459 3737
rect 3517 3737 3532 3743
rect 3485 3704 3491 3716
rect 3469 3584 3475 3696
rect 3469 3504 3475 3556
rect 3485 3544 3491 3696
rect 3501 3684 3507 3696
rect 3485 3484 3491 3536
rect 3453 3384 3459 3476
rect 3405 3317 3420 3323
rect 3389 3284 3395 3316
rect 3357 3044 3363 3056
rect 3293 2924 3299 2936
rect 3245 2777 3267 2783
rect 3108 2697 3123 2703
rect 3197 2644 3203 2696
rect 3112 2606 3118 2614
rect 3126 2606 3132 2614
rect 3140 2606 3146 2614
rect 3154 2606 3160 2614
rect 3181 2584 3187 2636
rect 3213 2584 3219 2696
rect 3229 2624 3235 2756
rect 3245 2704 3251 2716
rect 3261 2683 3267 2777
rect 3245 2677 3267 2683
rect 3117 2484 3123 2536
rect 3149 2524 3155 2576
rect 3172 2557 3196 2563
rect 3197 2524 3203 2556
rect 3213 2537 3228 2543
rect 3085 2304 3091 2316
rect 3005 2223 3011 2296
rect 2989 2217 3011 2223
rect 2989 2184 2995 2217
rect 2893 2044 2899 2096
rect 2909 2084 2915 2096
rect 2925 2084 2931 2116
rect 2941 2084 2947 2136
rect 2957 2103 2963 2156
rect 3005 2124 3011 2136
rect 2957 2097 2972 2103
rect 3005 2024 3011 2116
rect 3021 2024 3027 2276
rect 3037 2244 3043 2296
rect 3053 2264 3059 2276
rect 3069 2264 3075 2276
rect 3101 2264 3107 2416
rect 3117 2384 3123 2476
rect 3133 2364 3139 2496
rect 3165 2484 3171 2516
rect 3213 2484 3219 2537
rect 3245 2504 3251 2677
rect 3261 2604 3267 2636
rect 3293 2624 3299 2716
rect 3309 2684 3315 2936
rect 3357 2924 3363 2936
rect 3325 2684 3331 2916
rect 3341 2703 3347 2916
rect 3357 2744 3363 2776
rect 3341 2697 3356 2703
rect 3341 2644 3347 2676
rect 3373 2644 3379 3156
rect 3389 3024 3395 3216
rect 3421 3144 3427 3256
rect 3437 3204 3443 3316
rect 3453 3304 3459 3356
rect 3469 3164 3475 3336
rect 3501 3184 3507 3636
rect 3517 3484 3523 3737
rect 3741 3737 3756 3743
rect 3533 3704 3539 3716
rect 3421 3104 3427 3116
rect 3437 3104 3443 3116
rect 3469 3104 3475 3136
rect 3405 3097 3420 3103
rect 3405 3004 3411 3097
rect 3517 3103 3523 3316
rect 3533 3264 3539 3616
rect 3549 3504 3555 3696
rect 3565 3524 3571 3736
rect 3677 3704 3683 3716
rect 3581 3584 3587 3676
rect 3597 3524 3603 3536
rect 3565 3484 3571 3516
rect 3549 3303 3555 3456
rect 3613 3444 3619 3516
rect 3629 3504 3635 3576
rect 3549 3297 3571 3303
rect 3549 3184 3555 3276
rect 3565 3163 3571 3297
rect 3597 3284 3603 3436
rect 3629 3384 3635 3476
rect 3645 3424 3651 3496
rect 3677 3464 3683 3496
rect 3677 3384 3683 3416
rect 3629 3304 3635 3336
rect 3549 3157 3571 3163
rect 3517 3097 3532 3103
rect 3453 3064 3459 3076
rect 3421 2984 3427 2996
rect 3405 2964 3411 2976
rect 3437 2944 3443 3016
rect 3453 2924 3459 3016
rect 3389 2804 3395 2896
rect 3405 2844 3411 2916
rect 3469 2904 3475 3036
rect 3405 2723 3411 2836
rect 3396 2717 3411 2723
rect 3261 2544 3267 2576
rect 3149 2323 3155 2376
rect 3229 2324 3235 2476
rect 3261 2424 3267 2516
rect 3277 2364 3283 2616
rect 3309 2543 3315 2636
rect 3325 2623 3331 2636
rect 3325 2617 3356 2623
rect 3389 2584 3395 2676
rect 3309 2537 3347 2543
rect 3293 2424 3299 2496
rect 3309 2464 3315 2516
rect 3341 2484 3347 2537
rect 3325 2324 3331 2336
rect 3133 2317 3155 2323
rect 3133 2284 3139 2317
rect 3149 2244 3155 2296
rect 3165 2283 3171 2316
rect 3181 2304 3187 2316
rect 3165 2277 3187 2283
rect 3181 2263 3187 2277
rect 3181 2257 3196 2263
rect 3165 2243 3171 2256
rect 3165 2237 3187 2243
rect 3037 2224 3043 2236
rect 3037 2184 3043 2196
rect 3053 2144 3059 2156
rect 3037 1984 3043 2036
rect 3053 1984 3059 2136
rect 3069 2104 3075 2156
rect 3085 2084 3091 2236
rect 3181 2224 3187 2237
rect 3112 2206 3118 2214
rect 3126 2206 3132 2214
rect 3140 2206 3146 2214
rect 3154 2206 3160 2214
rect 3197 2124 3203 2256
rect 3213 2204 3219 2316
rect 3357 2304 3363 2556
rect 3373 2503 3379 2536
rect 3389 2524 3395 2536
rect 3405 2504 3411 2616
rect 3421 2563 3427 2876
rect 3437 2624 3443 2716
rect 3453 2663 3459 2896
rect 3469 2704 3475 2756
rect 3485 2744 3491 2896
rect 3501 2884 3507 3076
rect 3517 3064 3523 3076
rect 3533 3044 3539 3096
rect 3549 2964 3555 3157
rect 3581 3124 3587 3256
rect 3597 3144 3603 3276
rect 3565 3044 3571 3116
rect 3613 3063 3619 3276
rect 3645 3124 3651 3296
rect 3613 3057 3635 3063
rect 3517 2824 3523 2896
rect 3533 2804 3539 2896
rect 3549 2784 3555 2816
rect 3565 2764 3571 2876
rect 3581 2844 3587 2936
rect 3597 2924 3603 2976
rect 3613 2944 3619 3016
rect 3629 2804 3635 3057
rect 3581 2744 3587 2776
rect 3501 2717 3516 2723
rect 3453 2657 3475 2663
rect 3469 2644 3475 2657
rect 3453 2563 3459 2636
rect 3485 2563 3491 2716
rect 3501 2663 3507 2717
rect 3533 2684 3539 2716
rect 3501 2657 3523 2663
rect 3421 2557 3443 2563
rect 3453 2557 3475 2563
rect 3485 2557 3507 2563
rect 3437 2544 3443 2557
rect 3373 2497 3388 2503
rect 3261 2283 3267 2296
rect 3252 2277 3267 2283
rect 3229 2144 3235 2176
rect 3245 2144 3251 2256
rect 3293 2217 3308 2223
rect 3261 2184 3267 2216
rect 3181 2117 3196 2123
rect 3101 2044 3107 2116
rect 3133 2044 3139 2076
rect 2925 1924 2931 1956
rect 2845 1784 2851 1876
rect 2893 1804 2899 1876
rect 2813 1657 2835 1663
rect 2813 1644 2819 1657
rect 2813 1524 2819 1636
rect 2829 1544 2835 1636
rect 2845 1604 2851 1736
rect 2861 1684 2867 1716
rect 2861 1584 2867 1676
rect 2877 1604 2883 1796
rect 2941 1784 2947 1976
rect 3069 1943 3075 1976
rect 2996 1937 3011 1943
rect 2957 1924 2963 1936
rect 3005 1923 3011 1937
rect 3037 1937 3075 1943
rect 3005 1917 3027 1923
rect 3021 1884 3027 1917
rect 3037 1904 3043 1937
rect 2893 1524 2899 1536
rect 2909 1503 2915 1736
rect 2957 1723 2963 1796
rect 2973 1784 2979 1856
rect 2948 1717 2972 1723
rect 2925 1624 2931 1676
rect 2973 1664 2979 1696
rect 2893 1497 2915 1503
rect 2813 1444 2819 1496
rect 2877 1464 2883 1496
rect 2813 1324 2819 1396
rect 2845 1304 2851 1376
rect 2861 1344 2867 1436
rect 2877 1424 2883 1456
rect 2861 1324 2867 1336
rect 2797 1244 2803 1276
rect 2813 1264 2819 1296
rect 2813 1204 2819 1256
rect 2829 1204 2835 1296
rect 2877 1284 2883 1316
rect 2893 1304 2899 1497
rect 2925 1483 2931 1556
rect 2941 1524 2947 1616
rect 2989 1584 2995 1876
rect 3053 1864 3059 1916
rect 3053 1843 3059 1856
rect 3037 1837 3059 1843
rect 3005 1764 3011 1776
rect 3021 1704 3027 1796
rect 3037 1703 3043 1837
rect 3069 1824 3075 1896
rect 3085 1844 3091 1936
rect 3101 1924 3107 2016
rect 3149 1944 3155 2076
rect 3165 1984 3171 2036
rect 3181 1964 3187 2117
rect 3229 2064 3235 2096
rect 3197 2023 3203 2056
rect 3197 2017 3235 2023
rect 3117 1844 3123 1916
rect 3165 1904 3171 1936
rect 3053 1724 3059 1736
rect 3085 1723 3091 1836
rect 3112 1806 3118 1814
rect 3126 1806 3132 1814
rect 3140 1806 3146 1814
rect 3154 1806 3160 1814
rect 3085 1717 3100 1723
rect 3037 1697 3059 1703
rect 3053 1684 3059 1697
rect 3069 1584 3075 1696
rect 2957 1524 2963 1556
rect 3069 1544 3075 1556
rect 2973 1537 3059 1543
rect 2973 1503 2979 1537
rect 2964 1497 2979 1503
rect 3037 1484 3043 1516
rect 3053 1503 3059 1537
rect 3101 1524 3107 1676
rect 3053 1497 3084 1503
rect 3117 1503 3123 1776
rect 3181 1744 3187 1896
rect 3197 1884 3203 1956
rect 3213 1924 3219 1956
rect 3229 1864 3235 2017
rect 3261 1984 3267 2116
rect 3277 2064 3283 2196
rect 3293 2184 3299 2217
rect 3341 2144 3347 2296
rect 3373 2184 3379 2497
rect 3453 2464 3459 2536
rect 3469 2523 3475 2557
rect 3501 2524 3507 2557
rect 3469 2517 3491 2523
rect 3469 2464 3475 2496
rect 3485 2404 3491 2517
rect 3373 2144 3379 2156
rect 3341 2084 3347 2096
rect 3293 1943 3299 2076
rect 3325 1963 3331 2036
rect 3325 1957 3347 1963
rect 3277 1937 3299 1943
rect 3309 1937 3324 1943
rect 3261 1864 3267 1936
rect 3277 1904 3283 1937
rect 3197 1764 3203 1836
rect 3229 1784 3235 1856
rect 3277 1784 3283 1876
rect 3309 1864 3315 1937
rect 3341 1923 3347 1957
rect 3341 1917 3363 1923
rect 3357 1904 3363 1917
rect 3373 1884 3379 2136
rect 3389 2104 3395 2236
rect 3405 2184 3411 2376
rect 3453 2323 3459 2356
rect 3469 2343 3475 2396
rect 3485 2384 3491 2396
rect 3469 2337 3484 2343
rect 3453 2317 3468 2323
rect 3437 2284 3443 2316
rect 3453 2264 3459 2296
rect 3405 2144 3411 2156
rect 3437 2144 3443 2256
rect 3453 2144 3459 2156
rect 3469 2140 3475 2316
rect 3501 2304 3507 2476
rect 3517 2424 3523 2657
rect 3533 2544 3539 2596
rect 3549 2584 3555 2736
rect 3597 2664 3603 2776
rect 3645 2764 3651 2936
rect 3661 2743 3667 3376
rect 3709 3344 3715 3736
rect 3741 3584 3747 3737
rect 3773 3704 3779 3736
rect 3773 3604 3779 3696
rect 3741 3523 3747 3556
rect 3725 3517 3747 3523
rect 3725 3384 3731 3517
rect 3741 3444 3747 3496
rect 3757 3484 3763 3516
rect 3764 3477 3779 3483
rect 3773 3464 3779 3477
rect 3693 3304 3699 3336
rect 3725 3304 3731 3316
rect 3677 3284 3683 3296
rect 3725 3284 3731 3296
rect 3700 3077 3715 3083
rect 3709 2984 3715 3077
rect 3725 2904 3731 3276
rect 3741 3204 3747 3356
rect 3773 3324 3779 3396
rect 3805 3344 3811 4056
rect 3853 3924 3859 4096
rect 3853 3864 3859 3896
rect 3821 3824 3827 3856
rect 3821 3784 3827 3796
rect 3869 3756 3875 4136
rect 3885 3924 3891 3996
rect 3901 3904 3907 3916
rect 3917 3864 3923 3896
rect 3901 3784 3907 3816
rect 3933 3744 3939 4116
rect 3949 3924 3955 3956
rect 3965 3824 3971 4276
rect 4029 4184 4035 4317
rect 4077 4264 4083 4316
rect 4141 4264 4147 4496
rect 4157 4384 4163 4496
rect 4173 4484 4179 4516
rect 4189 4484 4195 4536
rect 4237 4484 4243 4516
rect 4253 4484 4259 4536
rect 4285 4464 4291 4496
rect 4189 4384 4195 4436
rect 4189 4337 4204 4343
rect 3981 4084 3987 4136
rect 3988 4077 4003 4083
rect 3981 3944 3987 3976
rect 3997 3904 4003 4077
rect 4077 4064 4083 4256
rect 4141 4184 4147 4236
rect 4109 4124 4115 4136
rect 4125 4104 4131 4156
rect 4173 4144 4179 4216
rect 4189 4184 4195 4337
rect 4205 4324 4211 4336
rect 4253 4284 4259 4316
rect 4301 4284 4307 4556
rect 4397 4544 4403 4636
rect 4413 4564 4419 4656
rect 4445 4624 4451 4896
rect 4477 4884 4483 5096
rect 4557 5064 4563 5116
rect 4573 5084 4579 5117
rect 4637 5104 4643 5117
rect 4717 5104 4723 5116
rect 4605 5084 4611 5096
rect 4621 5063 4627 5096
rect 4612 5057 4627 5063
rect 4573 5044 4579 5056
rect 4605 4984 4611 5056
rect 4733 5044 4739 5116
rect 4749 5104 4755 5136
rect 4765 5084 4771 5116
rect 4829 5104 4835 5136
rect 4845 5064 4851 5136
rect 4861 5084 4867 5257
rect 4893 5184 4899 5296
rect 4925 5224 4931 5316
rect 4957 5264 4963 5296
rect 4909 5144 4915 5156
rect 4797 5044 4803 5056
rect 4877 5044 4883 5116
rect 4941 5104 4947 5156
rect 4973 5104 4979 5316
rect 4989 5184 4995 5236
rect 5021 5224 5027 5296
rect 5053 5184 5059 5337
rect 5069 5324 5075 5336
rect 5085 5264 5091 5316
rect 5133 5304 5139 5496
rect 5165 5484 5171 5636
rect 5229 5544 5235 5756
rect 5405 5724 5411 5756
rect 5613 5724 5619 5843
rect 5629 5837 5651 5843
rect 5821 5837 5827 5843
rect 5869 5837 5875 5843
rect 5981 5837 6003 5843
rect 5629 5784 5635 5837
rect 5997 5764 6003 5837
rect 6093 5837 6115 5843
rect 5837 5744 5843 5756
rect 5917 5744 5923 5756
rect 5517 5704 5523 5716
rect 5613 5704 5619 5716
rect 5661 5683 5667 5716
rect 5661 5677 5676 5683
rect 5325 5504 5331 5576
rect 5405 5564 5411 5636
rect 5229 5464 5235 5476
rect 5341 5464 5347 5516
rect 5357 5464 5363 5536
rect 5389 5484 5395 5516
rect 5421 5464 5427 5576
rect 5437 5524 5443 5576
rect 5805 5564 5811 5718
rect 5901 5704 5907 5736
rect 5453 5504 5459 5536
rect 5469 5504 5475 5536
rect 5517 5524 5523 5536
rect 5549 5524 5555 5536
rect 5693 5524 5699 5536
rect 5789 5524 5795 5556
rect 5661 5517 5676 5523
rect 5181 5304 5187 5336
rect 5133 5264 5139 5276
rect 5149 5204 5155 5236
rect 5005 5104 5011 5116
rect 5021 5104 5027 5156
rect 4957 5084 4963 5096
rect 4941 4984 4947 5076
rect 5037 5064 5043 5136
rect 5037 5044 5043 5056
rect 5165 5043 5171 5276
rect 5213 5264 5219 5356
rect 5245 5284 5251 5456
rect 5533 5444 5539 5496
rect 5565 5444 5571 5516
rect 5597 5484 5603 5496
rect 5613 5464 5619 5476
rect 5405 5384 5411 5436
rect 5517 5424 5523 5436
rect 5661 5384 5667 5517
rect 5709 5504 5715 5516
rect 5837 5504 5843 5516
rect 5869 5504 5875 5696
rect 5933 5584 5939 5636
rect 5677 5484 5683 5496
rect 5725 5384 5731 5456
rect 5805 5424 5811 5476
rect 5901 5464 5907 5476
rect 5917 5464 5923 5496
rect 5917 5384 5923 5456
rect 5949 5364 5955 5456
rect 5981 5384 5987 5536
rect 5997 5384 6003 5496
rect 6045 5364 6051 5716
rect 6061 5584 6067 5696
rect 6061 5484 6067 5496
rect 5357 5304 5363 5356
rect 5469 5324 5475 5336
rect 5149 5037 5171 5043
rect 4989 4984 4995 5036
rect 5085 4984 5091 5036
rect 5149 4984 5155 5037
rect 5181 4984 5187 5216
rect 5245 5164 5251 5236
rect 5277 5124 5283 5296
rect 5341 5283 5347 5296
rect 5341 5277 5363 5283
rect 5341 5184 5347 5236
rect 5357 5144 5363 5277
rect 5437 5264 5443 5316
rect 5485 5304 5491 5316
rect 5485 5263 5491 5296
rect 5501 5264 5507 5296
rect 5533 5284 5539 5336
rect 5549 5304 5555 5316
rect 5581 5304 5587 5336
rect 5693 5324 5699 5336
rect 5709 5324 5715 5336
rect 5613 5304 5619 5316
rect 5469 5257 5491 5263
rect 5213 4984 5219 5096
rect 4541 4924 4547 4936
rect 4557 4904 4563 4976
rect 4573 4944 4579 4956
rect 4653 4944 4659 4956
rect 4861 4944 4867 4956
rect 4957 4944 4963 4976
rect 4733 4924 4739 4936
rect 4781 4904 4787 4916
rect 4605 4884 4611 4896
rect 4573 4784 4579 4836
rect 4632 4806 4638 4814
rect 4646 4806 4652 4814
rect 4660 4806 4666 4814
rect 4674 4806 4680 4814
rect 4829 4784 4835 4796
rect 4941 4784 4947 4936
rect 5021 4924 5027 4936
rect 4973 4904 4979 4916
rect 4989 4804 4995 4896
rect 5021 4784 5027 4916
rect 5037 4904 5043 4936
rect 5037 4864 5043 4896
rect 5085 4784 5091 4896
rect 4461 4704 4467 4716
rect 4477 4704 4483 4736
rect 4532 4717 4547 4723
rect 4493 4704 4499 4716
rect 4461 4584 4467 4656
rect 4509 4584 4515 4696
rect 4541 4604 4547 4717
rect 4573 4704 4579 4756
rect 4589 4584 4595 4716
rect 4605 4704 4611 4756
rect 4621 4684 4627 4736
rect 4637 4704 4643 4716
rect 4653 4664 4659 4676
rect 4605 4584 4611 4596
rect 4733 4584 4739 4676
rect 4765 4664 4771 4716
rect 4781 4704 4787 4716
rect 4797 4704 4803 4776
rect 4813 4684 4819 4736
rect 4845 4704 4851 4776
rect 5117 4744 5123 4916
rect 5165 4903 5171 4936
rect 5213 4904 5219 4916
rect 5156 4897 5171 4903
rect 5229 4903 5235 5036
rect 5245 4924 5251 5116
rect 5437 5104 5443 5176
rect 5453 5144 5459 5196
rect 5469 5184 5475 5257
rect 5565 5244 5571 5296
rect 5645 5263 5651 5316
rect 5741 5284 5747 5356
rect 5949 5344 5955 5356
rect 5789 5324 5795 5336
rect 5821 5324 5827 5336
rect 5885 5324 5891 5336
rect 5917 5324 5923 5336
rect 5757 5283 5763 5316
rect 5805 5284 5811 5296
rect 5821 5284 5827 5316
rect 5757 5277 5772 5283
rect 5741 5264 5747 5276
rect 5645 5257 5667 5263
rect 5485 5124 5491 5176
rect 5517 5144 5523 5196
rect 5501 5104 5507 5136
rect 5613 5124 5619 5256
rect 5629 5124 5635 5236
rect 5661 5184 5667 5257
rect 5757 5184 5763 5277
rect 5773 5184 5779 5256
rect 5853 5184 5859 5276
rect 5677 5144 5683 5156
rect 5741 5144 5747 5156
rect 5949 5124 5955 5316
rect 5981 5304 5987 5356
rect 5340 5064 5348 5070
rect 5261 5044 5267 5056
rect 5293 5044 5299 5056
rect 5229 4897 5244 4903
rect 5149 4784 5155 4876
rect 5197 4804 5203 4896
rect 5053 4737 5068 4743
rect 4765 4584 4771 4636
rect 4829 4584 4835 4656
rect 4893 4584 4899 4676
rect 4909 4624 4915 4696
rect 4989 4684 4995 4736
rect 5037 4684 5043 4696
rect 4925 4644 4931 4656
rect 4973 4584 4979 4616
rect 4989 4604 4995 4676
rect 5053 4664 5059 4737
rect 5076 4697 5084 4703
rect 5021 4624 5027 4636
rect 4349 4464 4355 4536
rect 4413 4524 4419 4556
rect 4493 4524 4499 4576
rect 4861 4544 4867 4556
rect 5005 4544 5011 4556
rect 5021 4544 5027 4556
rect 4541 4524 4547 4536
rect 4509 4464 4515 4496
rect 4253 4184 4259 4276
rect 4045 3964 4051 4036
rect 4093 3984 4099 4076
rect 4109 4064 4115 4096
rect 4125 4064 4131 4096
rect 4125 4004 4131 4056
rect 4141 3984 4147 4076
rect 4013 3924 4019 3956
rect 4045 3924 4051 3936
rect 4173 3924 4179 4096
rect 4205 3984 4211 4116
rect 4237 4103 4243 4156
rect 4237 4097 4252 4103
rect 4093 3904 4099 3916
rect 3981 3884 3987 3896
rect 4045 3784 4051 3876
rect 4157 3824 4163 3916
rect 4173 3904 4179 3916
rect 4189 3784 4195 3816
rect 4237 3784 4243 3896
rect 4285 3864 4291 4136
rect 4365 4103 4371 4156
rect 4356 4097 4371 4103
rect 4397 4084 4403 4136
rect 4413 4124 4419 4416
rect 4525 4384 4531 4436
rect 4541 4424 4547 4516
rect 4557 4464 4563 4536
rect 4701 4504 4707 4536
rect 4632 4406 4638 4414
rect 4646 4406 4652 4414
rect 4660 4406 4666 4414
rect 4674 4406 4680 4414
rect 4701 4384 4707 4496
rect 4749 4483 4755 4496
rect 4749 4477 4764 4483
rect 4765 4384 4771 4476
rect 4445 4263 4451 4316
rect 4429 4257 4451 4263
rect 4429 4184 4435 4257
rect 4477 4263 4483 4276
rect 4589 4264 4595 4276
rect 4477 4257 4499 4263
rect 4493 4184 4499 4257
rect 4557 4184 4563 4236
rect 4605 4184 4611 4256
rect 4685 4184 4691 4296
rect 4717 4283 4723 4316
rect 4717 4277 4732 4283
rect 4733 4204 4739 4276
rect 4484 4157 4499 4163
rect 4461 4144 4467 4156
rect 4301 3944 4307 3956
rect 4333 3944 4339 4036
rect 4397 3984 4403 4036
rect 4333 3904 4339 3916
rect 4349 3904 4355 3916
rect 4365 3884 4371 3956
rect 4429 3944 4435 4096
rect 4445 3984 4451 4116
rect 4461 3963 4467 4136
rect 4493 4104 4499 4157
rect 4525 4144 4531 4156
rect 4477 3984 4483 4076
rect 4461 3957 4483 3963
rect 4445 3904 4451 3956
rect 4477 3903 4483 3957
rect 4461 3897 4483 3903
rect 3837 3644 3843 3736
rect 3837 3584 3843 3596
rect 3933 3564 3939 3736
rect 3981 3704 3987 3736
rect 4013 3724 4019 3736
rect 4077 3724 4083 3756
rect 4157 3724 4163 3756
rect 3965 3697 3980 3703
rect 3965 3584 3971 3697
rect 3853 3464 3859 3476
rect 3869 3464 3875 3496
rect 3821 3324 3827 3396
rect 3837 3344 3843 3416
rect 3869 3384 3875 3436
rect 3901 3404 3907 3476
rect 3964 3464 3972 3470
rect 3997 3424 4003 3476
rect 4013 3444 4019 3716
rect 4061 3564 4067 3696
rect 4077 3664 4083 3696
rect 4157 3664 4163 3696
rect 4173 3564 4179 3696
rect 4189 3664 4195 3696
rect 4205 3644 4211 3676
rect 4237 3664 4243 3736
rect 4253 3724 4259 3736
rect 4205 3584 4211 3636
rect 4253 3584 4259 3716
rect 4301 3704 4307 3736
rect 4109 3464 4115 3476
rect 4125 3444 4131 3476
rect 4205 3404 4211 3496
rect 4045 3384 4051 3396
rect 4221 3384 4227 3476
rect 3853 3364 3859 3376
rect 3773 3204 3779 3316
rect 3741 3044 3747 3196
rect 3757 3124 3763 3156
rect 3789 3144 3795 3296
rect 3821 3184 3827 3316
rect 3885 3184 3891 3336
rect 3933 3324 3939 3356
rect 3981 3304 3987 3316
rect 3997 3304 4003 3316
rect 3965 3244 3971 3276
rect 3917 3224 3923 3236
rect 3853 3084 3859 3156
rect 3869 3124 3875 3176
rect 3885 3124 3891 3176
rect 3901 3124 3907 3196
rect 3917 3124 3923 3176
rect 3949 3164 3955 3236
rect 3981 3184 3987 3296
rect 4013 3244 4019 3316
rect 4029 3304 4035 3336
rect 4061 3324 4067 3356
rect 4221 3344 4227 3356
rect 4237 3324 4243 3476
rect 3901 3104 3907 3116
rect 3997 3104 4003 3116
rect 4013 3104 4019 3116
rect 4029 3104 4035 3136
rect 4061 3123 4067 3216
rect 4077 3204 4083 3296
rect 4093 3124 4099 3136
rect 4061 3117 4076 3123
rect 4029 3084 4035 3096
rect 3677 2763 3683 2856
rect 3677 2757 3699 2763
rect 3661 2737 3683 2743
rect 3645 2704 3651 2736
rect 3661 2664 3667 2716
rect 3613 2624 3619 2656
rect 3629 2584 3635 2656
rect 3556 2537 3580 2543
rect 3533 2524 3539 2536
rect 3597 2524 3603 2536
rect 3533 2484 3539 2496
rect 3517 2284 3523 2316
rect 3549 2264 3555 2496
rect 3581 2424 3587 2476
rect 3613 2464 3619 2576
rect 3581 2324 3587 2416
rect 3613 2344 3619 2376
rect 3629 2323 3635 2536
rect 3661 2464 3667 2536
rect 3677 2523 3683 2737
rect 3693 2544 3699 2757
rect 3725 2684 3731 2776
rect 3741 2764 3747 2936
rect 3709 2544 3715 2616
rect 3741 2584 3747 2696
rect 3757 2624 3763 3076
rect 3773 2764 3779 3056
rect 3789 2984 3795 3076
rect 3853 3064 3859 3076
rect 3869 3044 3875 3076
rect 3853 2944 3859 2996
rect 3869 2944 3875 2956
rect 3837 2924 3843 2936
rect 3837 2904 3843 2916
rect 3805 2744 3811 2856
rect 3837 2844 3843 2896
rect 3821 2744 3827 2756
rect 3869 2744 3875 2856
rect 3885 2784 3891 2836
rect 3837 2684 3843 2716
rect 3917 2704 3923 3036
rect 3949 3024 3955 3076
rect 3965 3064 3971 3076
rect 4061 3064 4067 3117
rect 4093 2984 4099 3076
rect 4109 3064 4115 3316
rect 4157 3144 4163 3156
rect 4173 3144 4179 3156
rect 4189 3124 4195 3236
rect 4237 3204 4243 3296
rect 4013 2924 4019 2976
rect 4029 2944 4035 2956
rect 4013 2884 4019 2916
rect 3933 2724 3939 2856
rect 3949 2784 3955 2836
rect 3965 2724 3971 2736
rect 3917 2664 3923 2676
rect 3725 2544 3731 2556
rect 3741 2524 3747 2536
rect 3757 2524 3763 2536
rect 3677 2517 3699 2523
rect 3629 2317 3651 2323
rect 3597 2284 3603 2316
rect 3437 1984 3443 2056
rect 3309 1784 3315 1856
rect 3277 1723 3283 1736
rect 3236 1717 3283 1723
rect 3197 1584 3203 1636
rect 3101 1497 3123 1503
rect 2916 1477 2931 1483
rect 3101 1483 3107 1497
rect 3133 1484 3139 1556
rect 3181 1517 3219 1523
rect 3149 1484 3155 1516
rect 3181 1503 3187 1517
rect 3165 1497 3187 1503
rect 3085 1477 3107 1483
rect 3005 1464 3011 1476
rect 2621 1084 2627 1096
rect 2765 1084 2771 1136
rect 2781 1064 2787 1116
rect 2845 1104 2851 1236
rect 2861 1164 2867 1236
rect 2925 1224 2931 1416
rect 2973 1404 2979 1436
rect 2957 1364 2963 1376
rect 2989 1324 2995 1456
rect 3005 1344 3011 1416
rect 3021 1324 3027 1476
rect 3085 1424 3091 1477
rect 3165 1464 3171 1497
rect 3213 1484 3219 1517
rect 3229 1484 3235 1616
rect 3277 1584 3283 1616
rect 3245 1544 3251 1576
rect 3261 1524 3267 1556
rect 3261 1504 3267 1516
rect 3112 1406 3118 1414
rect 3126 1406 3132 1414
rect 3140 1406 3146 1414
rect 3154 1406 3160 1414
rect 3181 1404 3187 1476
rect 3213 1444 3219 1476
rect 3085 1324 3091 1356
rect 2941 1244 2947 1316
rect 3197 1304 3203 1436
rect 3213 1304 3219 1336
rect 3245 1304 3251 1436
rect 3261 1384 3267 1496
rect 3293 1384 3299 1696
rect 3309 1504 3315 1556
rect 3325 1424 3331 1876
rect 3389 1864 3395 1916
rect 3373 1857 3388 1863
rect 3341 1824 3347 1836
rect 3357 1744 3363 1796
rect 3341 1724 3347 1736
rect 3373 1704 3379 1857
rect 3437 1784 3443 1896
rect 3453 1844 3459 1876
rect 3389 1584 3395 1736
rect 3341 1524 3347 1536
rect 3341 1484 3347 1516
rect 3373 1484 3379 1556
rect 3405 1424 3411 1676
rect 3453 1664 3459 1776
rect 3469 1543 3475 2076
rect 3485 1964 3491 2256
rect 3533 2164 3539 2176
rect 3501 1904 3507 1956
rect 3549 1904 3555 2236
rect 3565 2184 3571 2276
rect 3613 2264 3619 2276
rect 3533 1897 3548 1903
rect 3533 1864 3539 1897
rect 3549 1864 3555 1876
rect 3453 1537 3475 1543
rect 2877 1104 2883 1156
rect 2909 1104 2915 1136
rect 3021 1124 3027 1156
rect 3037 1123 3043 1276
rect 3277 1264 3283 1336
rect 3357 1324 3363 1376
rect 3165 1184 3171 1236
rect 3037 1117 3059 1123
rect 2797 1084 2803 1096
rect 2813 1063 2819 1096
rect 2893 1083 2899 1096
rect 2893 1077 2908 1083
rect 2925 1083 2931 1116
rect 2916 1077 2931 1083
rect 2797 1057 2819 1063
rect 2589 1004 2595 1056
rect 2797 1043 2803 1057
rect 2957 1044 2963 1116
rect 2973 1084 2979 1116
rect 3037 1044 3043 1056
rect 2612 1037 2803 1043
rect 2621 964 2627 976
rect 2589 904 2595 916
rect 2653 904 2659 916
rect 2564 877 2579 883
rect 2685 864 2691 896
rect 2701 863 2707 956
rect 2692 857 2707 863
rect 2484 717 2499 723
rect 2509 703 2515 716
rect 2500 697 2515 703
rect 2333 664 2339 676
rect 2381 624 2387 676
rect 2349 584 2355 596
rect 2397 564 2403 636
rect 2413 584 2419 656
rect 2461 644 2467 696
rect 2445 564 2451 636
rect 2477 584 2483 656
rect 2509 644 2515 676
rect 2541 664 2547 736
rect 2557 564 2563 656
rect 2237 504 2243 536
rect 2285 504 2291 536
rect 1901 304 1907 316
rect 1821 224 1827 296
rect 1837 184 1843 296
rect 1853 244 1859 276
rect 1933 264 1939 296
rect 1949 284 1955 356
rect 2237 344 2243 496
rect 2269 484 2275 496
rect 2381 484 2387 536
rect 2397 524 2403 536
rect 2429 504 2435 556
rect 2061 284 2067 316
rect 1853 184 1859 216
rect 1453 104 1459 116
rect 1853 104 1859 156
rect 1453 -17 1459 96
rect 1560 6 1566 14
rect 1574 6 1580 14
rect 1588 6 1594 14
rect 1602 6 1608 14
rect 1453 -23 1475 -17
rect 1869 -23 1875 256
rect 1981 144 1987 156
rect 2045 144 2051 156
rect 1965 -23 1971 96
rect 1981 -17 1987 136
rect 1997 104 2003 116
rect 2093 -17 2099 256
rect 2109 224 2115 276
rect 2141 204 2147 316
rect 2237 264 2243 296
rect 2285 264 2291 276
rect 2301 184 2307 436
rect 2349 184 2355 396
rect 2445 384 2451 536
rect 2509 524 2515 556
rect 2525 524 2531 536
rect 2509 484 2515 516
rect 2541 504 2547 556
rect 2573 544 2579 836
rect 2701 824 2707 857
rect 2717 764 2723 936
rect 2653 644 2659 696
rect 2669 684 2675 756
rect 2701 664 2707 736
rect 2669 604 2675 636
rect 2685 584 2691 616
rect 2733 584 2739 1016
rect 2909 984 2915 1016
rect 2989 984 2995 996
rect 2861 964 2867 976
rect 2829 924 2835 956
rect 3021 944 3027 996
rect 2861 924 2867 936
rect 2797 884 2803 916
rect 2781 864 2787 876
rect 2749 584 2755 796
rect 2765 784 2771 836
rect 2797 804 2803 876
rect 2845 744 2851 836
rect 2861 784 2867 896
rect 3053 884 3059 1117
rect 3069 1044 3075 1116
rect 3085 1104 3091 1176
rect 3101 1124 3107 1136
rect 3181 1084 3187 1236
rect 3293 1204 3299 1256
rect 3309 1184 3315 1296
rect 3341 1284 3347 1296
rect 3325 1184 3331 1196
rect 3197 1144 3203 1156
rect 3229 1124 3235 1176
rect 3357 1144 3363 1236
rect 3373 1224 3379 1396
rect 3405 1364 3411 1416
rect 3421 1404 3427 1436
rect 3421 1324 3427 1376
rect 3453 1364 3459 1537
rect 3485 1504 3491 1856
rect 3565 1783 3571 2076
rect 3581 2044 3587 2156
rect 3597 2144 3603 2156
rect 3597 2084 3603 2136
rect 3613 1964 3619 2176
rect 3645 2104 3651 2317
rect 3661 2204 3667 2316
rect 3677 2124 3683 2136
rect 3677 2084 3683 2096
rect 3636 2077 3660 2083
rect 3677 2064 3683 2076
rect 3629 1984 3635 2056
rect 3677 1964 3683 2036
rect 3581 1864 3587 1916
rect 3549 1777 3571 1783
rect 3501 1764 3507 1776
rect 3549 1724 3555 1777
rect 3549 1704 3555 1716
rect 3517 1424 3523 1476
rect 3533 1424 3539 1616
rect 3549 1524 3555 1616
rect 3581 1544 3587 1636
rect 3597 1484 3603 1776
rect 3613 1764 3619 1796
rect 3629 1764 3635 1896
rect 3661 1884 3667 1896
rect 3645 1804 3651 1876
rect 3613 1744 3619 1756
rect 3645 1704 3651 1756
rect 3613 1523 3619 1656
rect 3645 1524 3651 1636
rect 3613 1517 3635 1523
rect 3581 1444 3587 1476
rect 3613 1463 3619 1496
rect 3597 1457 3619 1463
rect 3485 1324 3491 1336
rect 3501 1303 3507 1376
rect 3533 1344 3539 1356
rect 3485 1297 3507 1303
rect 3469 1264 3475 1296
rect 3485 1263 3491 1297
rect 3485 1257 3507 1263
rect 3213 1104 3219 1116
rect 3245 1104 3251 1136
rect 3325 1124 3331 1136
rect 3373 1124 3379 1216
rect 3261 1084 3267 1116
rect 3325 1084 3331 1096
rect 3405 1084 3411 1136
rect 3485 1124 3491 1236
rect 3501 1123 3507 1257
rect 3517 1184 3523 1276
rect 3533 1124 3539 1216
rect 3549 1144 3555 1236
rect 3565 1184 3571 1436
rect 3581 1204 3587 1376
rect 3597 1344 3603 1457
rect 3629 1384 3635 1517
rect 3661 1503 3667 1776
rect 3677 1764 3683 1916
rect 3693 1784 3699 2517
rect 3725 2464 3731 2496
rect 3725 2424 3731 2456
rect 3725 2264 3731 2276
rect 3741 2244 3747 2456
rect 3773 2444 3779 2556
rect 3805 2464 3811 2536
rect 3821 2484 3827 2616
rect 3837 2544 3843 2656
rect 3933 2584 3939 2716
rect 3949 2684 3955 2716
rect 3981 2704 3987 2736
rect 4029 2724 4035 2936
rect 4093 2924 4099 2956
rect 4125 2940 4131 2996
rect 4061 2864 4067 2916
rect 4109 2903 4115 2936
rect 4100 2897 4115 2903
rect 4093 2744 4099 2896
rect 4045 2704 4051 2736
rect 3965 2664 3971 2696
rect 3981 2584 3987 2696
rect 4029 2664 4035 2696
rect 4077 2684 4083 2736
rect 4109 2684 4115 2716
rect 4125 2704 4131 2736
rect 3837 2504 3843 2536
rect 3885 2524 3891 2556
rect 3933 2544 3939 2556
rect 3901 2504 3907 2516
rect 3869 2464 3875 2476
rect 3885 2464 3891 2476
rect 3981 2444 3987 2516
rect 3997 2404 4003 2536
rect 4045 2504 4051 2636
rect 4061 2544 4067 2576
rect 4093 2564 4099 2636
rect 4077 2504 4083 2556
rect 3940 2337 3964 2343
rect 3757 2244 3763 2336
rect 3789 2224 3795 2316
rect 3837 2244 3843 2296
rect 3885 2264 3891 2316
rect 4013 2303 4019 2436
rect 4045 2304 4051 2396
rect 4068 2317 4083 2323
rect 3997 2297 4019 2303
rect 3917 2264 3923 2296
rect 3997 2244 4003 2297
rect 4029 2224 4035 2296
rect 4077 2284 4083 2317
rect 4093 2264 4099 2296
rect 4109 2184 4115 2656
rect 4141 2644 4147 3016
rect 4157 2984 4163 3116
rect 4189 3064 4195 3116
rect 4205 3104 4211 3156
rect 4253 3124 4259 3436
rect 4269 3364 4275 3516
rect 4285 3384 4291 3476
rect 4317 3384 4323 3876
rect 4333 3784 4339 3876
rect 4397 3864 4403 3896
rect 4397 3824 4403 3856
rect 4397 3784 4403 3796
rect 4429 3784 4435 3816
rect 4461 3784 4467 3897
rect 4493 3883 4499 4096
rect 4493 3877 4515 3883
rect 4493 3784 4499 3856
rect 4509 3784 4515 3877
rect 4525 3824 4531 3876
rect 4541 3804 4547 4096
rect 4557 3984 4563 4156
rect 4573 4144 4579 4176
rect 4829 4164 4835 4536
rect 4877 4504 4883 4516
rect 5053 4504 5059 4636
rect 5069 4584 5075 4696
rect 5101 4643 5107 4716
rect 5245 4704 5251 4716
rect 5117 4644 5123 4676
rect 5101 4637 5116 4643
rect 5213 4624 5219 4676
rect 5101 4584 5107 4596
rect 5085 4544 5091 4576
rect 5117 4564 5123 4576
rect 5229 4524 5235 4536
rect 4861 4184 4867 4496
rect 4973 4484 4979 4496
rect 5101 4384 5107 4496
rect 5133 4324 5139 4516
rect 5245 4344 5251 4536
rect 4877 4244 4883 4276
rect 4605 4104 4611 4116
rect 4589 3984 4595 4096
rect 4701 4084 4707 4156
rect 4893 4124 4899 4256
rect 4909 4124 4915 4136
rect 4925 4124 4931 4276
rect 4957 4263 4963 4316
rect 5117 4304 5123 4316
rect 4948 4257 4963 4263
rect 5005 4164 5011 4276
rect 4957 4124 4963 4136
rect 4632 4006 4638 4014
rect 4646 4006 4652 4014
rect 4660 4006 4666 4014
rect 4674 4006 4680 4014
rect 4701 3924 4707 4076
rect 4781 4044 4787 4116
rect 4845 4084 4851 4096
rect 4861 3944 4867 4096
rect 4893 3984 4899 4116
rect 4989 4104 4995 4116
rect 4941 4084 4947 4096
rect 4957 4064 4963 4076
rect 4909 3984 4915 4056
rect 4973 4044 4979 4096
rect 5005 4044 5011 4136
rect 5021 4064 5027 4296
rect 5101 4184 5107 4296
rect 5133 4284 5139 4316
rect 5037 4144 5043 4156
rect 5101 4124 5107 4136
rect 5005 3984 5011 4016
rect 5037 3984 5043 4116
rect 5053 4064 5059 4096
rect 5101 4024 5107 4116
rect 5117 4064 5123 4136
rect 5133 3984 5139 4256
rect 5165 4204 5171 4236
rect 5245 4224 5251 4236
rect 5229 4184 5235 4196
rect 5165 4144 5171 4176
rect 5245 4144 5251 4156
rect 5197 3964 5203 4116
rect 5245 4104 5251 4116
rect 5261 4064 5267 5016
rect 5341 4984 5347 5036
rect 5325 4944 5331 4956
rect 5277 4724 5283 4896
rect 5277 4584 5283 4716
rect 5309 4704 5315 4716
rect 5325 4664 5331 4936
rect 5405 4903 5411 5076
rect 5517 4984 5523 5116
rect 5549 4944 5555 5076
rect 5597 5063 5603 5076
rect 5629 5064 5635 5116
rect 5805 5084 5811 5096
rect 5821 5084 5827 5116
rect 5581 5057 5603 5063
rect 5581 4984 5587 5057
rect 5581 4964 5587 4976
rect 5437 4904 5443 4916
rect 5389 4897 5411 4903
rect 5341 4724 5347 4876
rect 5277 4504 5283 4536
rect 5277 4324 5283 4496
rect 5293 4384 5299 4656
rect 5341 4584 5347 4716
rect 5357 4504 5363 4616
rect 5373 4564 5379 4676
rect 5389 4384 5395 4897
rect 5405 4864 5411 4876
rect 5437 4844 5443 4896
rect 5453 4864 5459 4916
rect 5437 4784 5443 4816
rect 5485 4724 5491 4836
rect 5517 4684 5523 4736
rect 5533 4704 5539 4716
rect 5549 4704 5555 4936
rect 5581 4924 5587 4936
rect 5613 4924 5619 4956
rect 5565 4684 5571 4876
rect 5597 4824 5603 4896
rect 5629 4784 5635 5056
rect 5805 4984 5811 5076
rect 5741 4924 5747 4956
rect 5645 4744 5651 4876
rect 5661 4724 5667 4916
rect 5789 4884 5795 4956
rect 5485 4664 5491 4676
rect 5437 4584 5443 4636
rect 5581 4584 5587 4656
rect 5453 4544 5459 4556
rect 5428 4517 5443 4523
rect 5437 4384 5443 4517
rect 4573 3863 4579 3896
rect 4717 3884 4723 3916
rect 4893 3884 4899 3936
rect 4564 3857 4579 3863
rect 4557 3804 4563 3856
rect 4589 3763 4595 3856
rect 4605 3844 4611 3856
rect 4605 3784 4611 3796
rect 4637 3764 4643 3836
rect 4653 3824 4659 3876
rect 4717 3784 4723 3876
rect 4733 3784 4739 3836
rect 4589 3757 4611 3763
rect 4333 3724 4339 3736
rect 4413 3724 4419 3736
rect 4365 3644 4371 3716
rect 4452 3697 4467 3703
rect 4397 3584 4403 3696
rect 4461 3584 4467 3697
rect 4333 3524 4339 3576
rect 4445 3524 4451 3556
rect 4381 3464 4387 3516
rect 4493 3504 4499 3696
rect 4509 3584 4515 3756
rect 4541 3544 4547 3696
rect 4573 3564 4579 3716
rect 4589 3584 4595 3736
rect 4605 3584 4611 3757
rect 4637 3664 4643 3716
rect 4701 3624 4707 3776
rect 4749 3664 4755 3756
rect 4781 3724 4787 3796
rect 4632 3606 4638 3614
rect 4646 3606 4652 3614
rect 4660 3606 4666 3614
rect 4674 3606 4680 3614
rect 4397 3484 4403 3496
rect 4461 3484 4467 3496
rect 4381 3264 4387 3336
rect 4413 3104 4419 3396
rect 4461 3384 4467 3416
rect 4509 3384 4515 3476
rect 4685 3464 4691 3576
rect 4557 3404 4563 3456
rect 4621 3384 4627 3396
rect 4429 3284 4435 3296
rect 4429 3124 4435 3276
rect 4541 3164 4547 3336
rect 4557 3184 4563 3316
rect 4573 3297 4588 3303
rect 4573 3184 4579 3297
rect 4685 3284 4691 3456
rect 4221 3084 4227 3096
rect 4349 3044 4355 3076
rect 4237 2944 4243 3036
rect 4301 3004 4307 3036
rect 4189 2864 4195 2936
rect 4253 2924 4259 2996
rect 4285 2917 4300 2923
rect 4253 2884 4259 2916
rect 4173 2704 4179 2716
rect 4189 2704 4195 2856
rect 4253 2724 4259 2836
rect 4285 2744 4291 2917
rect 4397 2923 4403 3036
rect 4477 2984 4483 3096
rect 4525 3084 4531 3116
rect 4589 3104 4595 3276
rect 4632 3206 4638 3214
rect 4646 3206 4652 3214
rect 4660 3206 4666 3214
rect 4674 3206 4680 3214
rect 4701 3163 4707 3476
rect 4797 3384 4803 3776
rect 4829 3604 4835 3876
rect 4845 3764 4851 3816
rect 4909 3784 4915 3896
rect 4989 3784 4995 3936
rect 5005 3784 5011 3876
rect 5021 3864 5027 3916
rect 5085 3904 5091 3956
rect 4893 3704 4899 3756
rect 4909 3644 4915 3696
rect 4957 3584 4963 3716
rect 4813 3484 4819 3536
rect 4925 3524 4931 3536
rect 4893 3503 4899 3516
rect 4877 3497 4899 3503
rect 4877 3464 4883 3497
rect 4845 3424 4851 3456
rect 4829 3344 4835 3356
rect 4701 3157 4723 3163
rect 4388 2917 4403 2923
rect 4413 2884 4419 2896
rect 4429 2844 4435 2936
rect 4477 2904 4483 2956
rect 4381 2824 4387 2836
rect 4429 2784 4435 2836
rect 4301 2744 4307 2776
rect 4237 2704 4243 2716
rect 4285 2684 4291 2736
rect 4301 2704 4307 2716
rect 4317 2684 4323 2756
rect 4333 2704 4339 2776
rect 4445 2763 4451 2776
rect 4461 2764 4467 2896
rect 4477 2864 4483 2896
rect 4509 2884 4515 2936
rect 4477 2784 4483 2836
rect 4413 2757 4451 2763
rect 4413 2744 4419 2757
rect 4493 2744 4499 2836
rect 4525 2804 4531 3076
rect 4573 2984 4579 3056
rect 4589 3044 4595 3076
rect 4605 3064 4611 3136
rect 4621 3024 4627 3156
rect 4637 3064 4643 3096
rect 4701 3084 4707 3116
rect 4685 2944 4691 2976
rect 4701 2964 4707 3076
rect 4717 3063 4723 3157
rect 4829 3104 4835 3336
rect 4861 3184 4867 3336
rect 4797 3084 4803 3096
rect 4717 3057 4739 3063
rect 4717 2984 4723 3016
rect 4733 2984 4739 3057
rect 4749 3004 4755 3056
rect 4781 2984 4787 3076
rect 4541 2924 4547 2936
rect 4557 2924 4563 2936
rect 4781 2904 4787 2956
rect 4797 2924 4803 3076
rect 4813 2904 4819 2936
rect 4829 2904 4835 3056
rect 4861 3024 4867 3096
rect 4877 3064 4883 3356
rect 4893 3344 4899 3497
rect 4909 3424 4915 3496
rect 4925 3484 4931 3496
rect 4989 3384 4995 3476
rect 5005 3444 5011 3696
rect 5021 3684 5027 3856
rect 5053 3844 5059 3856
rect 5085 3784 5091 3896
rect 5133 3884 5139 3896
rect 5149 3884 5155 3896
rect 5245 3844 5251 3876
rect 5133 3784 5139 3836
rect 5053 3744 5059 3756
rect 5197 3744 5203 3836
rect 5277 3784 5283 4236
rect 5293 4184 5299 4296
rect 5325 4243 5331 4276
rect 5325 4237 5347 4243
rect 5309 4144 5315 4156
rect 5293 4024 5299 4096
rect 5309 3917 5324 3923
rect 5293 3844 5299 3876
rect 5309 3864 5315 3917
rect 5341 3883 5347 4237
rect 5405 4184 5411 4216
rect 5421 4184 5427 4276
rect 5405 4124 5411 4156
rect 5357 4084 5363 4096
rect 5405 4084 5411 4116
rect 5437 4064 5443 4336
rect 5453 4284 5459 4536
rect 5460 4257 5475 4263
rect 5325 3877 5347 3883
rect 5309 3784 5315 3856
rect 5325 3784 5331 3877
rect 5357 3844 5363 3876
rect 5373 3864 5379 3916
rect 5405 3863 5411 4056
rect 5469 3984 5475 4257
rect 5485 4084 5491 4576
rect 5565 4544 5571 4556
rect 5501 4517 5516 4523
rect 5501 4384 5507 4517
rect 5501 4124 5507 4296
rect 5517 4223 5523 4276
rect 5533 4244 5539 4396
rect 5549 4264 5555 4276
rect 5565 4243 5571 4516
rect 5597 4504 5603 4616
rect 5613 4584 5619 4676
rect 5661 4584 5667 4676
rect 5725 4664 5731 4876
rect 5805 4863 5811 4896
rect 5821 4884 5827 5076
rect 5869 4984 5875 5076
rect 5933 4964 5939 5116
rect 5981 5104 5987 5296
rect 6013 5184 6019 5316
rect 5949 5084 5955 5096
rect 5853 4884 5859 4936
rect 5885 4904 5891 4956
rect 5789 4857 5811 4863
rect 5741 4784 5747 4836
rect 5773 4764 5779 4816
rect 5789 4743 5795 4857
rect 5805 4764 5811 4836
rect 5853 4784 5859 4876
rect 5789 4737 5811 4743
rect 5741 4664 5747 4716
rect 5757 4704 5763 4736
rect 5805 4724 5811 4737
rect 5789 4704 5795 4716
rect 5677 4624 5683 4656
rect 5693 4584 5699 4656
rect 5709 4563 5715 4616
rect 5693 4557 5715 4563
rect 5581 4284 5587 4356
rect 5613 4344 5619 4536
rect 5613 4304 5619 4336
rect 5597 4297 5612 4303
rect 5581 4244 5587 4276
rect 5549 4237 5571 4243
rect 5517 4217 5539 4223
rect 5533 4164 5539 4217
rect 5501 3944 5507 4116
rect 5517 3884 5523 3916
rect 5533 3884 5539 4156
rect 5549 3883 5555 4237
rect 5597 4224 5603 4297
rect 5629 4284 5635 4296
rect 5693 4283 5699 4557
rect 5725 4524 5731 4536
rect 5677 4277 5699 4283
rect 5565 4184 5571 4196
rect 5629 4184 5635 4236
rect 5604 4117 5619 4123
rect 5581 3924 5587 3936
rect 5549 3877 5587 3883
rect 5389 3857 5411 3863
rect 5172 3717 5187 3723
rect 5085 3644 5091 3696
rect 5181 3664 5187 3717
rect 5245 3723 5251 3736
rect 5245 3717 5267 3723
rect 5117 3584 5123 3596
rect 5165 3584 5171 3656
rect 5197 3584 5203 3696
rect 5197 3524 5203 3536
rect 5085 3504 5091 3516
rect 5037 3384 5043 3496
rect 5053 3384 5059 3476
rect 5069 3424 5075 3456
rect 5117 3443 5123 3496
rect 5117 3437 5139 3443
rect 5005 3344 5011 3376
rect 4893 3304 4899 3316
rect 5021 3304 5027 3336
rect 5069 3323 5075 3336
rect 5117 3324 5123 3416
rect 5053 3317 5075 3323
rect 5053 3304 5059 3317
rect 4925 3184 4931 3256
rect 4989 3084 4995 3136
rect 4893 2984 4899 3076
rect 4925 2944 4931 2996
rect 4941 2984 4947 3036
rect 4957 2964 4963 2976
rect 4717 2884 4723 2896
rect 4509 2744 4515 2776
rect 4365 2704 4371 2716
rect 4349 2684 4355 2696
rect 4397 2684 4403 2716
rect 4429 2704 4435 2716
rect 4493 2704 4499 2736
rect 4509 2704 4515 2736
rect 4413 2684 4419 2696
rect 4141 2584 4147 2616
rect 4125 2384 4131 2436
rect 4141 2363 4147 2516
rect 4125 2357 4147 2363
rect 3741 2144 3747 2156
rect 3709 2044 3715 2096
rect 3741 2064 3747 2096
rect 3725 1904 3731 2016
rect 3709 1784 3715 1896
rect 3725 1864 3731 1876
rect 3677 1704 3683 1716
rect 3709 1704 3715 1756
rect 3725 1723 3731 1856
rect 3741 1744 3747 1896
rect 3725 1717 3740 1723
rect 3677 1564 3683 1636
rect 3661 1497 3683 1503
rect 3661 1464 3667 1476
rect 3613 1377 3628 1383
rect 3613 1344 3619 1377
rect 3629 1344 3635 1356
rect 3597 1324 3603 1336
rect 3645 1324 3651 1416
rect 3677 1383 3683 1497
rect 3661 1377 3683 1383
rect 3629 1317 3644 1323
rect 3597 1204 3603 1236
rect 3629 1203 3635 1317
rect 3661 1284 3667 1377
rect 3693 1363 3699 1496
rect 3741 1404 3747 1716
rect 3757 1583 3763 2176
rect 3821 2124 3827 2156
rect 3773 1724 3779 2096
rect 3789 2044 3795 2116
rect 3869 2084 3875 2156
rect 3901 2144 3907 2156
rect 3885 2137 3900 2143
rect 3885 2124 3891 2137
rect 3917 2124 3923 2176
rect 3965 2123 3971 2136
rect 3981 2124 3987 2156
rect 3949 2117 3971 2123
rect 3901 2103 3907 2116
rect 3949 2104 3955 2117
rect 3901 2097 3948 2103
rect 3821 1924 3827 1936
rect 3821 1784 3827 1836
rect 3869 1784 3875 1836
rect 3853 1724 3859 1776
rect 3901 1744 3907 2076
rect 3917 1984 3923 2036
rect 3940 1937 3955 1943
rect 3917 1824 3923 1896
rect 3933 1884 3939 1916
rect 3949 1904 3955 1937
rect 3997 1903 4003 2176
rect 4013 2104 4019 2116
rect 4029 1923 4035 2136
rect 4045 1964 4051 2116
rect 4125 2004 4131 2357
rect 4141 2284 4147 2316
rect 4141 2004 4147 2096
rect 4020 1917 4035 1923
rect 3997 1897 4019 1903
rect 3949 1864 3955 1896
rect 3965 1824 3971 1876
rect 3997 1864 4003 1876
rect 4013 1824 4019 1897
rect 4029 1884 4035 1917
rect 4061 1904 4067 1956
rect 4109 1903 4115 1976
rect 4109 1897 4124 1903
rect 4141 1903 4147 1996
rect 4157 1923 4163 2636
rect 4189 2584 4195 2596
rect 4205 2564 4211 2636
rect 4221 2404 4227 2596
rect 4429 2584 4435 2636
rect 4541 2584 4547 2876
rect 4589 2784 4595 2856
rect 4632 2806 4638 2814
rect 4646 2806 4652 2814
rect 4660 2806 4666 2814
rect 4674 2806 4680 2814
rect 4765 2804 4771 2896
rect 4829 2883 4835 2896
rect 4813 2877 4835 2883
rect 4573 2684 4579 2736
rect 4573 2644 4579 2676
rect 4653 2664 4659 2676
rect 4253 2524 4259 2536
rect 4253 2504 4259 2516
rect 4269 2504 4275 2556
rect 4397 2544 4403 2556
rect 4285 2504 4291 2536
rect 4333 2504 4339 2536
rect 4269 2464 4275 2496
rect 4317 2484 4323 2496
rect 4253 2404 4259 2436
rect 4173 2324 4179 2376
rect 4189 2284 4195 2316
rect 4205 2304 4211 2376
rect 4253 2324 4259 2396
rect 4285 2344 4291 2456
rect 4317 2264 4323 2416
rect 4381 2384 4387 2456
rect 4349 2304 4355 2316
rect 4365 2284 4371 2376
rect 4397 2284 4403 2476
rect 4413 2304 4419 2456
rect 4429 2324 4435 2496
rect 4445 2384 4451 2576
rect 4653 2544 4659 2556
rect 4557 2404 4563 2536
rect 4573 2504 4579 2516
rect 4573 2403 4579 2436
rect 4564 2397 4579 2403
rect 4589 2384 4595 2496
rect 4605 2424 4611 2536
rect 4685 2504 4691 2596
rect 4701 2564 4707 2696
rect 4765 2684 4771 2796
rect 4765 2663 4771 2676
rect 4756 2657 4771 2663
rect 4797 2663 4803 2696
rect 4813 2684 4819 2877
rect 4989 2844 4995 2956
rect 5021 2903 5027 3256
rect 5053 3104 5059 3296
rect 5101 3244 5107 3316
rect 5069 3064 5075 3196
rect 5069 2984 5075 3056
rect 5085 2924 5091 3216
rect 5117 3204 5123 3316
rect 5101 2944 5107 2976
rect 5005 2897 5027 2903
rect 5005 2884 5011 2897
rect 5021 2844 5027 2876
rect 4861 2724 4867 2776
rect 4845 2663 4851 2696
rect 4797 2657 4851 2663
rect 4632 2406 4638 2414
rect 4646 2406 4652 2414
rect 4660 2406 4666 2414
rect 4674 2406 4680 2414
rect 4701 2383 4707 2396
rect 4717 2384 4723 2596
rect 4740 2517 4764 2523
rect 4685 2377 4707 2383
rect 4605 2304 4611 2336
rect 4429 2284 4435 2296
rect 4653 2284 4659 2376
rect 4589 2264 4595 2276
rect 4173 2163 4179 2236
rect 4221 2204 4227 2256
rect 4461 2244 4467 2256
rect 4253 2237 4268 2243
rect 4237 2204 4243 2236
rect 4189 2163 4195 2176
rect 4221 2164 4227 2176
rect 4173 2157 4195 2163
rect 4173 2084 4179 2136
rect 4189 2124 4195 2157
rect 4253 2144 4259 2237
rect 4269 2144 4275 2216
rect 4397 2144 4403 2236
rect 4445 2184 4451 2196
rect 4509 2184 4515 2196
rect 4253 2124 4259 2136
rect 4269 2124 4275 2136
rect 4205 2104 4211 2116
rect 4285 2044 4291 2136
rect 4301 2124 4307 2136
rect 4413 2124 4419 2176
rect 4477 2124 4483 2176
rect 4301 2004 4307 2116
rect 4445 2104 4451 2116
rect 4509 2104 4515 2136
rect 4605 2124 4611 2136
rect 4669 2124 4675 2296
rect 4685 2184 4691 2377
rect 4733 2263 4739 2436
rect 4749 2363 4755 2436
rect 4765 2424 4771 2496
rect 4781 2384 4787 2636
rect 4877 2584 4883 2636
rect 4797 2484 4803 2556
rect 4813 2504 4819 2536
rect 4797 2363 4803 2476
rect 4813 2424 4819 2496
rect 4829 2484 4835 2536
rect 4845 2484 4851 2576
rect 4893 2563 4899 2756
rect 4909 2684 4915 2756
rect 4941 2644 4947 2836
rect 4973 2784 4979 2836
rect 5005 2784 5011 2836
rect 5053 2804 5059 2896
rect 5069 2884 5075 2896
rect 5005 2764 5011 2776
rect 5069 2764 5075 2876
rect 5101 2784 5107 2896
rect 5044 2717 5068 2723
rect 4973 2664 4979 2716
rect 5021 2584 5027 2696
rect 5053 2684 5059 2717
rect 5101 2703 5107 2756
rect 5085 2697 5107 2703
rect 5037 2644 5043 2676
rect 5085 2564 5091 2697
rect 4877 2557 4899 2563
rect 4877 2504 4883 2557
rect 4941 2524 4947 2536
rect 4829 2403 4835 2416
rect 4813 2397 4835 2403
rect 4813 2384 4819 2397
rect 4877 2384 4883 2496
rect 4925 2484 4931 2496
rect 4925 2457 4931 2476
rect 4941 2384 4947 2436
rect 4957 2384 4963 2476
rect 4749 2357 4803 2363
rect 4749 2304 4755 2316
rect 4765 2304 4771 2316
rect 4797 2297 4812 2303
rect 4717 2257 4739 2263
rect 4717 2224 4723 2257
rect 4733 2164 4739 2236
rect 4765 2224 4771 2276
rect 4781 2184 4787 2296
rect 4797 2244 4803 2297
rect 4829 2284 4835 2376
rect 4525 2104 4531 2116
rect 4381 2044 4387 2096
rect 4509 2084 4515 2096
rect 4541 2084 4547 2116
rect 4541 2064 4547 2076
rect 4557 2064 4563 2076
rect 4317 1944 4323 2036
rect 4349 1924 4355 2016
rect 4157 1917 4179 1923
rect 4173 1904 4179 1917
rect 4132 1897 4147 1903
rect 4125 1863 4131 1876
rect 4157 1864 4163 1896
rect 4116 1857 4131 1863
rect 4061 1784 4067 1816
rect 4141 1784 4147 1796
rect 3773 1604 3779 1716
rect 3757 1577 3779 1583
rect 3757 1504 3763 1556
rect 3773 1524 3779 1577
rect 3789 1524 3795 1656
rect 3805 1604 3811 1696
rect 3869 1684 3875 1736
rect 3933 1644 3939 1756
rect 4013 1744 4019 1756
rect 4061 1744 4067 1776
rect 3885 1624 3891 1636
rect 3949 1604 3955 1736
rect 3981 1703 3987 1716
rect 3981 1697 4003 1703
rect 3997 1644 4003 1697
rect 4077 1683 4083 1756
rect 4141 1744 4147 1776
rect 4109 1737 4124 1743
rect 4093 1684 4099 1696
rect 4077 1677 4092 1683
rect 4109 1644 4115 1737
rect 4125 1724 4131 1736
rect 4141 1683 4147 1716
rect 4157 1704 4163 1796
rect 4173 1743 4179 1896
rect 4189 1844 4195 1916
rect 4333 1904 4339 1916
rect 4221 1864 4227 1896
rect 4285 1844 4291 1856
rect 4365 1844 4371 1916
rect 4381 1904 4387 1916
rect 4397 1883 4403 2036
rect 4429 1884 4435 1916
rect 4445 1904 4451 1936
rect 4461 1884 4467 1896
rect 4381 1877 4403 1883
rect 4189 1744 4195 1796
rect 4173 1737 4188 1743
rect 4132 1677 4147 1683
rect 4125 1624 4131 1636
rect 3805 1584 3811 1596
rect 3853 1543 3859 1556
rect 3853 1537 3907 1543
rect 3805 1484 3811 1536
rect 3901 1524 3907 1537
rect 3901 1484 3907 1516
rect 3917 1484 3923 1576
rect 3933 1504 3939 1596
rect 3965 1524 3971 1616
rect 3949 1504 3955 1516
rect 3981 1484 3987 1596
rect 3677 1357 3699 1363
rect 3677 1324 3683 1357
rect 3709 1344 3715 1356
rect 3773 1344 3779 1376
rect 3789 1364 3795 1436
rect 3805 1384 3811 1436
rect 3869 1384 3875 1436
rect 3917 1364 3923 1416
rect 3693 1324 3699 1336
rect 3629 1197 3644 1203
rect 3501 1117 3516 1123
rect 3293 1064 3299 1076
rect 3325 1064 3331 1076
rect 3085 1037 3132 1043
rect 3085 1004 3091 1037
rect 3172 1037 3187 1043
rect 3181 1024 3187 1037
rect 3112 1006 3118 1014
rect 3126 1006 3132 1014
rect 3140 1006 3146 1014
rect 3154 1006 3160 1014
rect 3108 977 3219 983
rect 3117 944 3123 956
rect 3213 924 3219 977
rect 3229 924 3235 936
rect 3261 884 3267 996
rect 3277 984 3283 996
rect 3293 924 3299 936
rect 3293 904 3299 916
rect 2925 784 2931 856
rect 2765 724 2771 736
rect 2813 684 2819 736
rect 2845 684 2851 716
rect 2877 684 2883 696
rect 2909 684 2915 736
rect 2941 724 2947 876
rect 2957 704 2963 816
rect 3037 764 3043 876
rect 3021 717 3075 723
rect 3021 704 3027 717
rect 3069 704 3075 717
rect 2957 684 2963 696
rect 2973 684 2979 696
rect 2973 664 2979 676
rect 3021 664 3027 676
rect 3069 664 3075 676
rect 2765 584 2771 636
rect 2525 464 2531 496
rect 2541 424 2547 496
rect 2621 464 2627 536
rect 2717 484 2723 536
rect 2733 464 2739 536
rect 2797 524 2803 596
rect 2765 484 2771 496
rect 2813 444 2819 636
rect 2877 544 2883 556
rect 2877 524 2883 536
rect 2893 524 2899 596
rect 2941 524 2947 536
rect 3005 524 3011 536
rect 3021 524 3027 536
rect 2893 384 2899 456
rect 2957 384 2963 476
rect 3005 404 3011 516
rect 3069 504 3075 516
rect 2717 324 2723 336
rect 2413 164 2419 216
rect 1981 -23 2003 -17
rect 2077 -23 2099 -17
rect 2157 -23 2163 16
rect 2221 -17 2227 156
rect 2333 144 2339 156
rect 2381 144 2387 156
rect 2445 140 2451 236
rect 2237 124 2243 136
rect 2349 104 2355 116
rect 2205 -23 2227 -17
rect 2333 -23 2339 16
rect 2461 -23 2467 276
rect 2477 264 2483 316
rect 2493 184 2499 316
rect 2637 264 2643 316
rect 2797 284 2803 336
rect 2813 304 2819 316
rect 2749 264 2755 276
rect 2845 264 2851 336
rect 2909 284 2915 336
rect 2925 243 2931 276
rect 3069 264 3075 316
rect 3053 257 3068 263
rect 3037 244 3043 256
rect 2925 237 2947 243
rect 2829 224 2835 236
rect 2765 184 2771 196
rect 2941 184 2947 237
rect 2989 184 2995 236
rect 3053 184 3059 257
rect 3085 204 3091 816
rect 3181 624 3187 836
rect 3197 684 3203 736
rect 3213 704 3219 796
rect 3309 744 3315 776
rect 3197 664 3203 676
rect 3277 644 3283 716
rect 3341 704 3347 776
rect 3357 724 3363 1076
rect 3389 984 3395 1056
rect 3421 1044 3427 1076
rect 3437 1044 3443 1096
rect 3453 1004 3459 1076
rect 3469 1043 3475 1116
rect 3485 1084 3491 1116
rect 3533 1084 3539 1116
rect 3565 1103 3571 1156
rect 3597 1104 3603 1116
rect 3556 1097 3571 1103
rect 3613 1084 3619 1156
rect 3629 1063 3635 1156
rect 3661 1124 3667 1236
rect 3709 1184 3715 1276
rect 3789 1244 3795 1336
rect 3821 1284 3827 1296
rect 3757 1204 3763 1236
rect 3869 1224 3875 1316
rect 3885 1304 3891 1316
rect 3741 1144 3747 1196
rect 3661 1104 3667 1116
rect 3757 1104 3763 1156
rect 3645 1084 3651 1096
rect 3677 1077 3740 1083
rect 3565 1057 3635 1063
rect 3469 1037 3491 1043
rect 3485 1024 3491 1037
rect 3373 944 3379 956
rect 3389 824 3395 956
rect 3437 944 3443 956
rect 3469 924 3475 1016
rect 3549 964 3555 1036
rect 3565 1024 3571 1057
rect 3677 1063 3683 1077
rect 3652 1057 3683 1063
rect 3517 924 3523 936
rect 3581 924 3587 1016
rect 3773 984 3779 1116
rect 3805 1077 3820 1083
rect 3709 944 3715 956
rect 3805 944 3811 1077
rect 3828 1057 3859 1063
rect 3853 1024 3859 1057
rect 3837 984 3843 1016
rect 3869 984 3875 1036
rect 3885 1024 3891 1296
rect 3901 1284 3907 1316
rect 3901 1184 3907 1236
rect 3917 1224 3923 1336
rect 3917 1063 3923 1176
rect 3933 1143 3939 1416
rect 3949 1324 3955 1356
rect 3981 1343 3987 1376
rect 3972 1337 3987 1343
rect 3997 1324 4003 1496
rect 4045 1464 4051 1516
rect 4077 1364 4083 1596
rect 4093 1544 4099 1556
rect 4125 1524 4131 1536
rect 4173 1524 4179 1556
rect 4189 1484 4195 1736
rect 4205 1664 4211 1736
rect 4221 1724 4227 1816
rect 4317 1744 4323 1776
rect 4365 1744 4371 1796
rect 4221 1504 4227 1556
rect 4237 1524 4243 1716
rect 4269 1684 4275 1696
rect 4253 1504 4259 1576
rect 4269 1564 4275 1676
rect 4285 1504 4291 1516
rect 4285 1464 4291 1476
rect 3997 1164 4003 1316
rect 4013 1184 4019 1336
rect 4029 1304 4035 1316
rect 4045 1203 4051 1336
rect 4036 1197 4051 1203
rect 3933 1137 3955 1143
rect 3949 1124 3955 1137
rect 4029 1124 4035 1196
rect 4061 1123 4067 1356
rect 4077 1144 4083 1356
rect 4157 1344 4163 1396
rect 4173 1344 4179 1436
rect 4109 1324 4115 1336
rect 4189 1284 4195 1436
rect 4285 1424 4291 1436
rect 4205 1384 4211 1396
rect 4205 1304 4211 1316
rect 4269 1303 4275 1356
rect 4260 1297 4275 1303
rect 4125 1123 4131 1236
rect 4205 1224 4211 1296
rect 4301 1264 4307 1696
rect 4365 1504 4371 1576
rect 4317 1384 4323 1476
rect 4333 1384 4339 1436
rect 4349 1424 4355 1476
rect 4356 1417 4371 1423
rect 4365 1364 4371 1417
rect 4173 1184 4179 1216
rect 4205 1184 4211 1196
rect 4253 1124 4259 1256
rect 4349 1144 4355 1236
rect 4365 1184 4371 1236
rect 4381 1224 4387 1877
rect 4477 1864 4483 1916
rect 4557 1884 4563 1916
rect 4509 1864 4515 1876
rect 4541 1864 4547 1876
rect 4397 1744 4403 1796
rect 4461 1784 4467 1836
rect 4413 1684 4419 1696
rect 4397 1524 4403 1556
rect 4413 1524 4419 1676
rect 4429 1644 4435 1756
rect 4477 1744 4483 1756
rect 4525 1744 4531 1836
rect 4573 1804 4579 2116
rect 4589 2084 4595 2096
rect 4621 2064 4627 2076
rect 4632 2006 4638 2014
rect 4646 2006 4652 2014
rect 4660 2006 4666 2014
rect 4674 2006 4680 2014
rect 4701 1983 4707 2116
rect 4717 2044 4723 2156
rect 4733 2023 4739 2136
rect 4813 2124 4819 2276
rect 4829 2144 4835 2256
rect 4845 2164 4851 2276
rect 4941 2244 4947 2276
rect 4957 2264 4963 2316
rect 4765 2024 4771 2036
rect 4685 1977 4707 1983
rect 4717 2017 4739 2023
rect 4605 1904 4611 1956
rect 4621 1884 4627 1916
rect 4589 1844 4595 1876
rect 4653 1844 4659 1876
rect 4573 1784 4579 1796
rect 4573 1757 4588 1763
rect 4413 1444 4419 1456
rect 4397 1164 4403 1436
rect 4429 1324 4435 1576
rect 4461 1564 4467 1636
rect 4477 1604 4483 1716
rect 4573 1704 4579 1757
rect 4621 1743 4627 1836
rect 4612 1737 4627 1743
rect 4589 1724 4595 1736
rect 4685 1724 4691 1977
rect 4717 1704 4723 2017
rect 4829 2004 4835 2136
rect 4845 1964 4851 2136
rect 4893 2104 4899 2216
rect 4877 2083 4883 2096
rect 4861 2077 4883 2083
rect 4788 1937 4812 1943
rect 4845 1924 4851 1956
rect 4829 1904 4835 1916
rect 4749 1844 4755 1880
rect 4733 1724 4739 1756
rect 4765 1724 4771 1776
rect 4445 1324 4451 1356
rect 4420 1317 4428 1323
rect 4477 1264 4483 1596
rect 4509 1484 4515 1516
rect 4541 1504 4547 1656
rect 4557 1584 4563 1636
rect 4632 1606 4638 1614
rect 4646 1606 4652 1614
rect 4660 1606 4666 1614
rect 4674 1606 4680 1614
rect 4525 1464 4531 1496
rect 4557 1444 4563 1516
rect 4589 1504 4595 1516
rect 4589 1464 4595 1496
rect 4653 1484 4659 1576
rect 4717 1484 4723 1516
rect 4733 1504 4739 1696
rect 4749 1664 4755 1696
rect 4781 1684 4787 1856
rect 4813 1784 4819 1896
rect 4861 1884 4867 2077
rect 4877 1904 4883 1956
rect 4909 1924 4915 2236
rect 4957 2224 4963 2236
rect 4973 2203 4979 2476
rect 4989 2384 4995 2516
rect 5021 2303 5027 2396
rect 5037 2344 5043 2536
rect 5053 2464 5059 2556
rect 5085 2324 5091 2556
rect 5101 2484 5107 2656
rect 5117 2644 5123 3176
rect 5133 3124 5139 3437
rect 5149 3364 5155 3476
rect 5165 3424 5171 3496
rect 5197 3484 5203 3516
rect 5245 3504 5251 3516
rect 5261 3484 5267 3717
rect 5341 3584 5347 3616
rect 5357 3604 5363 3736
rect 5389 3644 5395 3857
rect 5421 3843 5427 3876
rect 5533 3864 5539 3876
rect 5421 3837 5443 3843
rect 5437 3784 5443 3837
rect 5501 3784 5507 3816
rect 5453 3684 5459 3736
rect 5277 3504 5283 3536
rect 5245 3464 5251 3476
rect 5213 3384 5219 3456
rect 5261 3364 5267 3476
rect 5293 3464 5299 3476
rect 5309 3463 5315 3496
rect 5309 3457 5324 3463
rect 5133 3104 5139 3116
rect 5133 2944 5139 2996
rect 5149 2924 5155 3356
rect 5181 3244 5187 3316
rect 5213 3284 5219 3296
rect 5165 3104 5171 3116
rect 5229 3104 5235 3316
rect 5293 3304 5299 3316
rect 5165 3084 5171 3096
rect 5181 3044 5187 3076
rect 5213 2964 5219 3056
rect 5229 2983 5235 3096
rect 5245 3084 5251 3236
rect 5261 3184 5267 3236
rect 5293 3164 5299 3296
rect 5309 3004 5315 3457
rect 5373 3444 5379 3496
rect 5325 3384 5331 3436
rect 5389 3384 5395 3476
rect 5405 3384 5411 3416
rect 5341 3304 5347 3356
rect 5357 3344 5363 3356
rect 5421 3224 5427 3636
rect 5437 3584 5443 3676
rect 5485 3644 5491 3736
rect 5517 3624 5523 3776
rect 5549 3744 5555 3756
rect 5533 3644 5539 3716
rect 5437 3464 5443 3496
rect 5453 3484 5459 3536
rect 5469 3464 5475 3516
rect 5325 3104 5331 3116
rect 5437 3084 5443 3316
rect 5453 3304 5459 3316
rect 5469 3184 5475 3296
rect 5229 2977 5251 2983
rect 5165 2924 5171 2936
rect 5197 2784 5203 2816
rect 5213 2784 5219 2816
rect 5133 2744 5139 2756
rect 5181 2723 5187 2776
rect 5197 2744 5203 2756
rect 5213 2723 5219 2756
rect 5181 2717 5219 2723
rect 5149 2624 5155 2696
rect 5133 2524 5139 2536
rect 5117 2464 5123 2496
rect 5021 2297 5043 2303
rect 4989 2264 4995 2280
rect 5021 2264 5027 2276
rect 4957 2197 4979 2203
rect 4941 2144 4947 2156
rect 4957 2123 4963 2197
rect 4973 2124 4979 2156
rect 4948 2117 4963 2123
rect 4925 1924 4931 2036
rect 4941 2004 4947 2116
rect 4989 2084 4995 2176
rect 5021 2124 5027 2176
rect 5037 2164 5043 2297
rect 5101 2263 5107 2316
rect 5117 2284 5123 2396
rect 5133 2304 5139 2516
rect 5165 2504 5171 2596
rect 5181 2344 5187 2636
rect 5213 2624 5219 2696
rect 5229 2564 5235 2956
rect 5245 2924 5251 2977
rect 5373 2944 5379 2976
rect 5405 2904 5411 3016
rect 5437 2984 5443 3076
rect 5453 2984 5459 3076
rect 5245 2797 5299 2803
rect 5245 2764 5251 2797
rect 5277 2744 5283 2776
rect 5293 2763 5299 2797
rect 5357 2784 5363 2836
rect 5389 2824 5395 2896
rect 5405 2824 5411 2896
rect 5421 2884 5427 2896
rect 5293 2757 5331 2763
rect 5252 2737 5267 2743
rect 5245 2664 5251 2716
rect 5261 2584 5267 2737
rect 5293 2704 5299 2736
rect 5309 2644 5315 2736
rect 5325 2723 5331 2757
rect 5325 2717 5372 2723
rect 5380 2717 5395 2723
rect 5348 2697 5372 2703
rect 5389 2684 5395 2717
rect 5437 2664 5443 2676
rect 5293 2564 5299 2596
rect 5213 2544 5219 2556
rect 5261 2537 5276 2543
rect 5245 2524 5251 2536
rect 5261 2503 5267 2537
rect 5204 2497 5267 2503
rect 5277 2484 5283 2496
rect 5277 2344 5283 2376
rect 5213 2324 5219 2336
rect 5309 2284 5315 2556
rect 5373 2544 5379 2556
rect 5325 2524 5331 2536
rect 5405 2503 5411 2596
rect 5437 2564 5443 2636
rect 5421 2504 5427 2536
rect 5437 2524 5443 2536
rect 5389 2497 5411 2503
rect 5389 2384 5395 2497
rect 5453 2384 5459 2936
rect 5469 2864 5475 2956
rect 5485 2784 5491 3616
rect 5565 3484 5571 3736
rect 5581 3724 5587 3877
rect 5597 3784 5603 4096
rect 5613 3984 5619 4117
rect 5629 4104 5635 4156
rect 5645 4124 5651 4236
rect 5661 4104 5667 4236
rect 5677 4164 5683 4277
rect 5709 4224 5715 4436
rect 5725 4324 5731 4496
rect 5741 4484 5747 4536
rect 5789 4524 5795 4596
rect 5805 4544 5811 4716
rect 5821 4544 5827 4736
rect 5853 4704 5859 4756
rect 5853 4604 5859 4696
rect 5869 4544 5875 4836
rect 5901 4784 5907 4916
rect 5933 4803 5939 4896
rect 5949 4864 5955 5076
rect 6045 4984 6051 5076
rect 6061 5064 6067 5356
rect 6093 5084 6099 5837
rect 6141 5784 6147 5843
rect 6173 5764 6179 5843
rect 6125 5684 6131 5696
rect 6141 5584 6147 5756
rect 6205 5717 6220 5723
rect 6173 5704 6179 5716
rect 6189 5684 6195 5696
rect 6109 5384 6115 5496
rect 6189 5324 6195 5436
rect 6205 5384 6211 5717
rect 6221 5364 6227 5636
rect 6237 5544 6243 5736
rect 6237 5323 6243 5496
rect 6221 5317 6243 5323
rect 6189 5224 6195 5296
rect 6205 5144 6211 5236
rect 6221 5184 6227 5317
rect 6253 5244 6259 5476
rect 6205 5063 6211 5116
rect 6189 5057 6211 5063
rect 6077 5044 6083 5056
rect 5965 4924 5971 4956
rect 5917 4797 5939 4803
rect 5885 4644 5891 4676
rect 5901 4664 5907 4716
rect 5917 4683 5923 4797
rect 5933 4704 5939 4756
rect 5949 4724 5955 4736
rect 5917 4677 5939 4683
rect 5901 4604 5907 4656
rect 5901 4584 5907 4596
rect 5933 4584 5939 4677
rect 5965 4624 5971 4896
rect 5981 4804 5987 4916
rect 5997 4884 6003 4976
rect 6029 4944 6035 4956
rect 6061 4923 6067 5036
rect 6109 4984 6115 4996
rect 6125 4956 6131 5036
rect 6189 4923 6195 5057
rect 6221 5003 6227 5056
rect 6237 5024 6243 5136
rect 6221 4997 6243 5003
rect 6045 4917 6067 4923
rect 6173 4917 6195 4923
rect 5981 4704 5987 4716
rect 5997 4643 6003 4856
rect 6045 4844 6051 4917
rect 6061 4844 6067 4896
rect 6061 4804 6067 4836
rect 6141 4784 6147 4836
rect 6045 4704 6051 4716
rect 6013 4664 6019 4696
rect 6061 4684 6067 4756
rect 5997 4637 6019 4643
rect 5981 4584 5987 4636
rect 5789 4484 5795 4496
rect 5805 4337 5820 4343
rect 5725 4304 5731 4316
rect 5805 4304 5811 4337
rect 5837 4304 5843 4536
rect 5885 4504 5891 4536
rect 5901 4504 5907 4576
rect 5917 4524 5923 4536
rect 5869 4497 5884 4503
rect 5741 4264 5747 4296
rect 5853 4284 5859 4476
rect 5869 4384 5875 4497
rect 5917 4364 5923 4516
rect 5933 4484 5939 4496
rect 5725 4164 5731 4236
rect 5677 4064 5683 4116
rect 5693 4104 5699 4156
rect 5709 4124 5715 4136
rect 5693 4023 5699 4076
rect 5725 4064 5731 4136
rect 5741 4103 5747 4216
rect 5741 4097 5763 4103
rect 5677 4017 5699 4023
rect 5613 3864 5619 3896
rect 5629 3744 5635 3876
rect 5661 3804 5667 3896
rect 5677 3784 5683 4017
rect 5693 3864 5699 3916
rect 5725 3824 5731 3876
rect 5693 3784 5699 3796
rect 5533 3344 5539 3436
rect 5581 3404 5587 3716
rect 5597 3583 5603 3736
rect 5613 3723 5619 3736
rect 5613 3717 5635 3723
rect 5613 3604 5619 3696
rect 5629 3664 5635 3717
rect 5645 3704 5651 3716
rect 5661 3683 5667 3776
rect 5741 3764 5747 3876
rect 5645 3677 5667 3683
rect 5597 3577 5619 3583
rect 5613 3344 5619 3577
rect 5645 3503 5651 3677
rect 5661 3524 5667 3556
rect 5645 3497 5667 3503
rect 5629 3384 5635 3396
rect 5645 3384 5651 3436
rect 5661 3364 5667 3497
rect 5517 3204 5523 3336
rect 5581 3324 5587 3336
rect 5549 3184 5555 3196
rect 5501 3104 5507 3116
rect 5501 3023 5507 3076
rect 5517 3044 5523 3076
rect 5501 3017 5523 3023
rect 5517 2984 5523 3017
rect 5533 2964 5539 3116
rect 5565 3064 5571 3076
rect 5533 2784 5539 2936
rect 5549 2924 5555 2956
rect 5565 2944 5571 3056
rect 5581 3024 5587 3296
rect 5597 3104 5603 3316
rect 5613 3104 5619 3156
rect 5629 3104 5635 3356
rect 5645 3184 5651 3316
rect 5661 3204 5667 3316
rect 5677 3264 5683 3656
rect 5725 3544 5731 3576
rect 5741 3564 5747 3756
rect 5757 3744 5763 4097
rect 5773 4004 5779 4236
rect 5789 4224 5795 4264
rect 5837 4184 5843 4256
rect 5853 4244 5859 4256
rect 5805 4104 5811 4136
rect 5821 4124 5827 4176
rect 5837 4104 5843 4136
rect 5869 4123 5875 4296
rect 5885 4284 5891 4296
rect 5917 4264 5923 4296
rect 5949 4264 5955 4316
rect 5901 4224 5907 4236
rect 5853 4117 5875 4123
rect 5773 3804 5779 3856
rect 5789 3724 5795 4096
rect 5805 3944 5811 3976
rect 5821 3904 5827 3996
rect 5837 3924 5843 3936
rect 5853 3883 5859 4117
rect 5869 4064 5875 4096
rect 5885 4084 5891 4116
rect 5869 4044 5875 4056
rect 5885 4004 5891 4036
rect 5901 4024 5907 4076
rect 5869 3944 5875 3976
rect 5901 3943 5907 3996
rect 5917 3964 5923 4036
rect 5933 4004 5939 4256
rect 5949 4244 5955 4256
rect 5965 4184 5971 4536
rect 5981 4484 5987 4536
rect 6013 4364 6019 4637
rect 5965 4064 5971 4116
rect 5901 3937 5923 3943
rect 5837 3877 5859 3883
rect 5821 3824 5827 3836
rect 5805 3744 5811 3756
rect 5821 3744 5827 3796
rect 5789 3604 5795 3676
rect 5773 3584 5779 3596
rect 5700 3477 5715 3483
rect 5709 3463 5715 3477
rect 5709 3457 5724 3463
rect 5693 3384 5699 3456
rect 5709 3384 5715 3457
rect 5741 3424 5747 3516
rect 5757 3464 5763 3536
rect 5789 3524 5795 3576
rect 5757 3404 5763 3456
rect 5773 3344 5779 3476
rect 5789 3424 5795 3456
rect 5709 3184 5715 3336
rect 5757 3284 5763 3336
rect 5789 3264 5795 3316
rect 5613 3084 5619 3096
rect 5597 3003 5603 3016
rect 5581 2997 5603 3003
rect 5549 2824 5555 2916
rect 5581 2903 5587 2997
rect 5629 2984 5635 3076
rect 5645 2984 5651 3136
rect 5661 3124 5667 3136
rect 5677 3104 5683 3116
rect 5661 2964 5667 3096
rect 5693 3064 5699 3116
rect 5709 3063 5715 3156
rect 5741 3124 5747 3236
rect 5805 3223 5811 3696
rect 5821 3664 5827 3716
rect 5837 3643 5843 3877
rect 5901 3864 5907 3916
rect 5853 3784 5859 3856
rect 5885 3783 5891 3836
rect 5917 3784 5923 3937
rect 5933 3864 5939 3936
rect 5949 3864 5955 3996
rect 5965 3904 5971 4036
rect 5981 4004 5987 4356
rect 6013 4304 6019 4316
rect 6013 4144 6019 4276
rect 6029 4264 6035 4656
rect 6045 4284 6051 4616
rect 6077 4564 6083 4716
rect 6157 4704 6163 4736
rect 6093 4604 6099 4656
rect 6093 4543 6099 4556
rect 6084 4537 6099 4543
rect 6061 4344 6067 4536
rect 6109 4524 6115 4696
rect 6173 4684 6179 4917
rect 6205 4884 6211 4916
rect 6141 4677 6156 4683
rect 6045 4224 6051 4256
rect 6077 4223 6083 4516
rect 6093 4504 6099 4516
rect 6125 4504 6131 4676
rect 6141 4564 6147 4677
rect 6189 4683 6195 4836
rect 6205 4704 6211 4836
rect 6221 4824 6227 4876
rect 6189 4677 6204 4683
rect 6157 4484 6163 4656
rect 6173 4544 6179 4656
rect 6109 4284 6115 4336
rect 6061 4217 6083 4223
rect 6045 4144 6051 4156
rect 6004 4097 6019 4103
rect 5981 3944 5987 3956
rect 5965 3884 5971 3896
rect 5885 3777 5907 3783
rect 5885 3724 5891 3756
rect 5853 3664 5859 3696
rect 5901 3683 5907 3777
rect 5933 3724 5939 3796
rect 5949 3764 5955 3836
rect 5965 3804 5971 3836
rect 5981 3804 5987 3856
rect 5965 3704 5971 3776
rect 5949 3684 5955 3696
rect 5901 3677 5916 3683
rect 5837 3637 5859 3643
rect 5837 3584 5843 3596
rect 5853 3543 5859 3637
rect 5997 3643 6003 4056
rect 6013 3844 6019 4097
rect 6061 4064 6067 4217
rect 6093 4104 6099 4256
rect 6125 4164 6131 4476
rect 6173 4424 6179 4496
rect 6141 4304 6147 4316
rect 6157 4284 6163 4376
rect 6189 4364 6195 4436
rect 6205 4324 6211 4356
rect 6221 4304 6227 4696
rect 6237 4624 6243 4997
rect 6253 4984 6259 5216
rect 6253 4904 6259 4936
rect 6253 4444 6259 4876
rect 6253 4284 6259 4396
rect 6109 4124 6115 4156
rect 6029 3984 6035 4036
rect 6077 3964 6083 4036
rect 6029 3944 6035 3956
rect 6061 3897 6076 3903
rect 6045 3884 6051 3896
rect 6029 3763 6035 3856
rect 6045 3783 6051 3836
rect 6061 3783 6067 3897
rect 6077 3824 6083 3876
rect 6045 3777 6067 3783
rect 6020 3757 6035 3763
rect 5981 3637 6003 3643
rect 5869 3584 5875 3636
rect 5853 3537 5875 3543
rect 5821 3497 5836 3503
rect 5821 3383 5827 3497
rect 5837 3404 5843 3456
rect 5853 3444 5859 3516
rect 5821 3377 5843 3383
rect 5821 3264 5827 3296
rect 5789 3217 5811 3223
rect 5725 3083 5731 3096
rect 5725 3077 5747 3083
rect 5709 3057 5731 3063
rect 5725 2963 5731 3057
rect 5741 2983 5747 3077
rect 5757 3064 5763 3116
rect 5773 3084 5779 3096
rect 5789 3024 5795 3217
rect 5837 3223 5843 3377
rect 5828 3217 5843 3223
rect 5821 3184 5827 3216
rect 5837 3184 5843 3196
rect 5821 3104 5827 3176
rect 5869 3144 5875 3537
rect 5885 3424 5891 3536
rect 5901 3344 5907 3496
rect 5917 3364 5923 3596
rect 5949 3484 5955 3576
rect 5981 3564 5987 3637
rect 5997 3584 6003 3616
rect 6013 3604 6019 3736
rect 6029 3684 6035 3757
rect 5933 3363 5939 3476
rect 5949 3444 5955 3456
rect 5949 3384 5955 3436
rect 5933 3357 5955 3363
rect 5885 3284 5891 3336
rect 5933 3304 5939 3336
rect 5949 3323 5955 3357
rect 5965 3344 5971 3556
rect 6045 3544 6051 3756
rect 6061 3724 6067 3777
rect 6077 3684 6083 3816
rect 5997 3504 6003 3536
rect 6061 3464 6067 3476
rect 6077 3444 6083 3656
rect 6093 3644 6099 4056
rect 6109 4024 6115 4096
rect 6141 4063 6147 4276
rect 6157 4244 6163 4276
rect 6189 4204 6195 4236
rect 6157 4157 6172 4163
rect 6157 4144 6163 4157
rect 6180 4137 6195 4143
rect 6141 4057 6156 4063
rect 6125 3984 6131 3996
rect 6141 3984 6147 4016
rect 6141 3864 6147 3956
rect 6157 3884 6163 4056
rect 6173 3964 6179 4096
rect 6189 4064 6195 4137
rect 6157 3844 6163 3856
rect 6109 3764 6115 3836
rect 6157 3803 6163 3836
rect 6141 3797 6163 3803
rect 6125 3784 6131 3796
rect 6141 3764 6147 3797
rect 6157 3744 6163 3776
rect 6109 3704 6115 3736
rect 6125 3664 6131 3716
rect 6141 3644 6147 3736
rect 6173 3704 6179 3856
rect 6189 3804 6195 4036
rect 6189 3744 6195 3776
rect 6109 3524 6115 3616
rect 6125 3504 6131 3636
rect 6141 3504 6147 3576
rect 6173 3524 6179 3696
rect 6189 3544 6195 3636
rect 6189 3484 6195 3496
rect 5981 3324 5987 3436
rect 5949 3317 5971 3323
rect 5917 3284 5923 3296
rect 5901 3264 5907 3276
rect 5885 3257 5900 3263
rect 5805 3084 5811 3096
rect 5837 3083 5843 3136
rect 5885 3124 5891 3257
rect 5901 3124 5907 3236
rect 5917 3184 5923 3216
rect 5869 3104 5875 3116
rect 5828 3077 5843 3083
rect 5757 3003 5763 3016
rect 5757 2997 5779 3003
rect 5741 2977 5763 2983
rect 5757 2964 5763 2977
rect 5725 2957 5740 2963
rect 5572 2897 5587 2903
rect 5581 2763 5587 2836
rect 5597 2824 5603 2936
rect 5613 2844 5619 2936
rect 5645 2923 5651 2956
rect 5773 2944 5779 2997
rect 5805 2984 5811 3056
rect 5837 3044 5843 3077
rect 5837 3024 5843 3036
rect 5805 2964 5811 2976
rect 5789 2943 5795 2956
rect 5789 2937 5811 2943
rect 5677 2924 5683 2936
rect 5725 2924 5731 2936
rect 5645 2917 5667 2923
rect 5661 2904 5667 2917
rect 5645 2883 5651 2896
rect 5645 2877 5683 2883
rect 5677 2864 5683 2877
rect 5533 2757 5587 2763
rect 5469 2724 5475 2756
rect 5501 2744 5507 2756
rect 5533 2743 5539 2757
rect 5517 2737 5539 2743
rect 5517 2703 5523 2737
rect 5492 2697 5523 2703
rect 5533 2684 5539 2716
rect 5661 2704 5667 2716
rect 5645 2664 5651 2696
rect 5613 2643 5619 2656
rect 5677 2644 5683 2856
rect 5693 2784 5699 2876
rect 5709 2743 5715 2896
rect 5725 2844 5731 2916
rect 5741 2784 5747 2936
rect 5805 2924 5811 2937
rect 5789 2904 5795 2916
rect 5757 2844 5763 2896
rect 5757 2824 5763 2836
rect 5805 2824 5811 2896
rect 5757 2784 5763 2816
rect 5773 2763 5779 2816
rect 5821 2784 5827 2976
rect 5869 2964 5875 2976
rect 5885 2943 5891 3036
rect 5869 2937 5891 2943
rect 5757 2757 5779 2763
rect 5757 2744 5763 2757
rect 5693 2737 5715 2743
rect 5693 2704 5699 2737
rect 5725 2704 5731 2716
rect 5741 2664 5747 2736
rect 5773 2724 5779 2736
rect 5757 2664 5763 2696
rect 5604 2637 5619 2643
rect 5469 2484 5475 2496
rect 5325 2324 5331 2336
rect 5437 2284 5443 2296
rect 5469 2284 5475 2316
rect 5277 2264 5283 2276
rect 5101 2257 5116 2263
rect 5053 2163 5059 2236
rect 5069 2184 5075 2236
rect 5053 2157 5068 2163
rect 5037 2144 5043 2156
rect 5053 2124 5059 2157
rect 5085 2124 5091 2256
rect 5325 2244 5331 2276
rect 5101 2144 5107 2176
rect 5133 2124 5139 2156
rect 5149 2144 5155 2196
rect 5213 2184 5219 2196
rect 5165 2123 5171 2156
rect 5245 2124 5251 2216
rect 5325 2144 5331 2176
rect 5293 2124 5299 2136
rect 5341 2124 5347 2156
rect 5389 2144 5395 2176
rect 5485 2164 5491 2636
rect 5549 2584 5555 2616
rect 5565 2577 5651 2583
rect 5565 2544 5571 2577
rect 5645 2556 5651 2577
rect 5597 2524 5603 2536
rect 5533 2504 5539 2516
rect 5517 2464 5523 2476
rect 5533 2424 5539 2496
rect 5549 2464 5555 2496
rect 5661 2484 5667 2516
rect 5581 2343 5587 2416
rect 5572 2337 5587 2343
rect 5581 2304 5587 2337
rect 5725 2323 5731 2636
rect 5741 2584 5747 2656
rect 5789 2624 5795 2776
rect 5837 2724 5843 2916
rect 5853 2844 5859 2936
rect 5869 2864 5875 2937
rect 5805 2584 5811 2716
rect 5789 2544 5795 2556
rect 5773 2497 5788 2503
rect 5773 2464 5779 2497
rect 5725 2317 5747 2323
rect 5549 2264 5555 2296
rect 5597 2264 5603 2276
rect 5629 2264 5635 2316
rect 5693 2284 5699 2316
rect 5645 2224 5651 2276
rect 5709 2224 5715 2276
rect 5741 2224 5747 2317
rect 5773 2283 5779 2316
rect 5789 2304 5795 2456
rect 5821 2384 5827 2676
rect 5853 2664 5859 2816
rect 5869 2744 5875 2836
rect 5901 2724 5907 2836
rect 5917 2743 5923 3156
rect 5933 2984 5939 3296
rect 5965 3283 5971 3317
rect 5997 3284 6003 3376
rect 5965 3277 5987 3283
rect 5981 3263 5987 3277
rect 6013 3263 6019 3276
rect 5981 3257 6019 3263
rect 5965 3184 5971 3256
rect 5949 2984 5955 3076
rect 5981 2964 5987 3156
rect 6013 3144 6019 3176
rect 6029 3124 6035 3416
rect 6061 3384 6067 3396
rect 6141 3364 6147 3396
rect 6173 3364 6179 3476
rect 6189 3343 6195 3456
rect 6205 3404 6211 4176
rect 6221 4084 6227 4096
rect 6237 4004 6243 4236
rect 6221 3784 6227 3896
rect 6237 3744 6243 3876
rect 6221 3664 6227 3696
rect 6221 3544 6227 3596
rect 6221 3384 6227 3456
rect 6173 3337 6195 3343
rect 6125 3324 6131 3336
rect 5997 3043 6003 3116
rect 6061 3044 6067 3276
rect 6077 3104 6083 3116
rect 5997 3037 6019 3043
rect 6013 2984 6019 3037
rect 5949 2924 5955 2956
rect 5981 2903 5987 2936
rect 5997 2904 6003 2976
rect 6013 2904 6019 2936
rect 5933 2897 5987 2903
rect 5933 2784 5939 2897
rect 5949 2824 5955 2876
rect 5917 2737 5939 2743
rect 5908 2717 5923 2723
rect 5837 2644 5843 2656
rect 5853 2624 5859 2636
rect 5885 2623 5891 2676
rect 5917 2664 5923 2717
rect 5885 2617 5916 2623
rect 5837 2603 5843 2616
rect 5837 2597 5875 2603
rect 5837 2544 5843 2556
rect 5853 2544 5859 2556
rect 5805 2344 5811 2356
rect 5773 2277 5795 2283
rect 5156 2117 5171 2123
rect 5005 2104 5011 2116
rect 5149 2084 5155 2116
rect 5277 2084 5283 2116
rect 5309 2084 5315 2096
rect 5357 2044 5363 2136
rect 5405 2124 5411 2156
rect 5389 2104 5395 2116
rect 5373 2044 5379 2096
rect 4989 2024 4995 2036
rect 4941 1903 4947 1956
rect 4957 1904 4963 2016
rect 5204 1917 5219 1923
rect 5149 1904 5155 1916
rect 4932 1897 4947 1903
rect 4861 1864 4867 1876
rect 4941 1804 4947 1876
rect 5037 1864 5043 1876
rect 4829 1744 4835 1796
rect 4989 1784 4995 1856
rect 5069 1764 5075 1836
rect 5133 1784 5139 1896
rect 5149 1864 5155 1876
rect 5213 1844 5219 1917
rect 5229 1864 5235 1876
rect 5213 1784 5219 1836
rect 5261 1764 5267 1976
rect 5373 1964 5379 2036
rect 5421 1964 5427 2116
rect 5437 2104 5443 2116
rect 5485 2084 5491 2116
rect 5517 2104 5523 2116
rect 5469 2044 5475 2076
rect 5485 2064 5491 2076
rect 5501 2044 5507 2096
rect 5533 2044 5539 2116
rect 5581 2084 5587 2136
rect 5613 2064 5619 2096
rect 5645 2064 5651 2216
rect 5757 2204 5763 2236
rect 5789 2184 5795 2277
rect 5661 2124 5667 2136
rect 5677 2104 5683 2116
rect 5773 2104 5779 2136
rect 5709 2084 5715 2096
rect 5725 2064 5731 2076
rect 5277 1864 5283 1876
rect 5293 1844 5299 1856
rect 5325 1844 5331 1896
rect 5373 1824 5379 1896
rect 5421 1884 5427 1956
rect 5453 1924 5459 2036
rect 5501 2024 5507 2036
rect 5469 1944 5475 1956
rect 5453 1903 5459 1916
rect 5485 1904 5491 1916
rect 5444 1897 5459 1903
rect 5533 1884 5539 2016
rect 5549 1924 5555 1936
rect 5533 1864 5539 1876
rect 5277 1784 5283 1816
rect 5549 1784 5555 1916
rect 5597 1903 5603 2036
rect 5629 1904 5635 2036
rect 5741 2024 5747 2096
rect 5805 2044 5811 2236
rect 5773 1984 5779 2016
rect 5677 1977 5731 1983
rect 5661 1904 5667 1916
rect 5597 1897 5619 1903
rect 5597 1864 5603 1876
rect 4973 1744 4979 1756
rect 5261 1744 5267 1756
rect 5293 1744 5299 1756
rect 4877 1737 4915 1743
rect 4813 1604 4819 1636
rect 4829 1564 4835 1736
rect 4877 1724 4883 1737
rect 4909 1723 4915 1737
rect 4909 1717 4931 1723
rect 4749 1484 4755 1496
rect 4637 1464 4643 1480
rect 4765 1464 4771 1516
rect 4861 1504 4867 1536
rect 4797 1444 4803 1476
rect 4845 1444 4851 1496
rect 4781 1424 4787 1436
rect 4493 1344 4499 1356
rect 4541 1344 4547 1416
rect 4541 1303 4547 1316
rect 4541 1297 4588 1303
rect 4525 1284 4531 1296
rect 4381 1124 4387 1136
rect 4061 1117 4083 1123
rect 4125 1117 4147 1123
rect 3997 1064 4003 1096
rect 4061 1064 4067 1096
rect 4077 1084 4083 1117
rect 4116 1097 4131 1103
rect 4077 1064 4083 1076
rect 3908 1057 3923 1063
rect 3821 964 3827 976
rect 3405 824 3411 896
rect 3357 684 3363 696
rect 3389 684 3395 756
rect 3437 724 3443 896
rect 3501 864 3507 896
rect 3453 703 3459 836
rect 3501 724 3507 736
rect 3437 697 3459 703
rect 3389 644 3395 656
rect 3112 606 3118 614
rect 3126 606 3132 614
rect 3140 606 3146 614
rect 3154 606 3160 614
rect 3149 484 3155 576
rect 3165 504 3171 516
rect 3181 504 3187 536
rect 3197 483 3203 516
rect 3213 504 3219 536
rect 3188 477 3203 483
rect 3165 464 3171 476
rect 3261 464 3267 536
rect 3293 524 3299 636
rect 3405 544 3411 616
rect 3437 584 3443 697
rect 3613 684 3619 916
rect 3677 904 3683 936
rect 3645 724 3651 896
rect 3725 744 3731 756
rect 3645 704 3651 716
rect 3773 684 3779 696
rect 3453 664 3459 676
rect 3421 544 3427 556
rect 3309 464 3315 536
rect 3421 324 3427 336
rect 3181 244 3187 296
rect 3325 284 3331 316
rect 3453 304 3459 656
rect 3485 344 3491 676
rect 3501 564 3507 636
rect 3581 584 3587 636
rect 3709 584 3715 616
rect 3789 584 3795 836
rect 3805 784 3811 816
rect 3837 764 3843 836
rect 3821 664 3827 696
rect 3853 664 3859 676
rect 3501 544 3507 556
rect 3613 544 3619 556
rect 3709 544 3715 556
rect 3725 544 3731 556
rect 3517 504 3523 536
rect 3693 444 3699 516
rect 3805 504 3811 536
rect 3837 524 3843 556
rect 3885 544 3891 1016
rect 3917 963 3923 1036
rect 4029 984 4035 1036
rect 4093 964 4099 1076
rect 4125 964 4131 1097
rect 3901 957 3923 963
rect 3901 904 3907 957
rect 3949 904 3955 956
rect 4093 924 4099 956
rect 4013 917 4028 923
rect 4013 904 4019 917
rect 3901 724 3907 756
rect 3917 724 3923 736
rect 3933 644 3939 856
rect 3949 684 3955 696
rect 3965 684 3971 736
rect 3997 704 4003 836
rect 4141 703 4147 1117
rect 4157 1083 4163 1096
rect 4157 1077 4179 1083
rect 4157 1004 4163 1056
rect 4173 943 4179 1077
rect 4189 1064 4195 1116
rect 4253 1064 4259 1096
rect 4413 1084 4419 1096
rect 4429 1063 4435 1116
rect 4413 1057 4435 1063
rect 4301 984 4307 1036
rect 4413 1024 4419 1057
rect 4365 984 4371 1016
rect 4429 964 4435 1036
rect 4445 984 4451 1236
rect 4493 1084 4499 1116
rect 4477 1044 4483 1076
rect 4605 1004 4611 1336
rect 4637 1304 4643 1336
rect 4717 1284 4723 1316
rect 4813 1303 4819 1356
rect 4804 1297 4819 1303
rect 4632 1206 4638 1214
rect 4646 1206 4652 1214
rect 4660 1206 4666 1214
rect 4674 1206 4680 1214
rect 4813 1184 4819 1297
rect 4861 1184 4867 1496
rect 4893 1484 4899 1716
rect 4925 1703 4931 1717
rect 5005 1703 5011 1716
rect 5037 1704 5043 1716
rect 4925 1697 5011 1703
rect 5085 1664 5091 1736
rect 5133 1704 5139 1736
rect 4957 1584 4963 1656
rect 5149 1624 5155 1736
rect 5357 1704 5363 1756
rect 5389 1724 5395 1736
rect 5261 1624 5267 1696
rect 5405 1684 5411 1716
rect 5485 1704 5491 1756
rect 5501 1724 5507 1736
rect 5597 1724 5603 1756
rect 5453 1644 5459 1676
rect 5469 1624 5475 1636
rect 5485 1603 5491 1696
rect 5469 1597 5491 1603
rect 4941 1504 4947 1516
rect 4957 1504 4963 1536
rect 4973 1484 4979 1516
rect 5005 1464 5011 1496
rect 5021 1464 5027 1516
rect 4877 1344 4883 1356
rect 5037 1344 5043 1596
rect 5469 1584 5475 1597
rect 5053 1344 5059 1456
rect 5085 1424 5091 1476
rect 5165 1464 5171 1516
rect 5309 1504 5315 1556
rect 5181 1424 5187 1476
rect 5325 1464 5331 1516
rect 5341 1504 5347 1536
rect 5357 1524 5363 1556
rect 5357 1484 5363 1516
rect 5405 1464 5411 1476
rect 5133 1340 5139 1396
rect 5245 1344 5251 1436
rect 5277 1384 5283 1456
rect 5421 1444 5427 1476
rect 5005 1324 5011 1336
rect 5268 1337 5292 1343
rect 5053 1264 5059 1316
rect 5101 1244 5107 1316
rect 4637 1104 4643 1116
rect 4781 1104 4787 1116
rect 4829 1084 4835 1116
rect 4749 1044 4755 1076
rect 4845 1064 4851 1096
rect 4925 1084 4931 1236
rect 4941 1084 4947 1156
rect 4957 1104 4963 1116
rect 4861 1044 4867 1076
rect 4973 1064 4979 1236
rect 4989 1064 4995 1156
rect 5053 1104 5059 1236
rect 5101 1084 5107 1236
rect 5149 1184 5155 1336
rect 5309 1324 5315 1436
rect 5421 1364 5427 1436
rect 5437 1384 5443 1496
rect 5469 1444 5475 1496
rect 5165 1304 5171 1316
rect 5245 1244 5251 1296
rect 5293 1244 5299 1316
rect 5421 1304 5427 1356
rect 5469 1344 5475 1436
rect 5437 1324 5443 1336
rect 5533 1304 5539 1476
rect 5581 1464 5587 1476
rect 5613 1464 5619 1897
rect 5677 1883 5683 1977
rect 5709 1904 5715 1956
rect 5725 1943 5731 1977
rect 5725 1937 5756 1943
rect 5725 1904 5731 1916
rect 5773 1884 5779 1896
rect 5668 1877 5683 1883
rect 5789 1844 5795 1916
rect 5821 1864 5827 2216
rect 5837 2183 5843 2516
rect 5869 2364 5875 2597
rect 5933 2563 5939 2737
rect 5949 2664 5955 2736
rect 5949 2604 5955 2656
rect 5981 2584 5987 2836
rect 6013 2764 6019 2896
rect 6013 2724 6019 2736
rect 6029 2704 6035 3036
rect 6061 2944 6067 3016
rect 6093 2984 6099 3096
rect 6125 3023 6131 3216
rect 6157 3124 6163 3236
rect 6157 3064 6163 3076
rect 6173 3064 6179 3337
rect 6237 3324 6243 3716
rect 6196 3137 6211 3143
rect 6205 3104 6211 3137
rect 6237 3124 6243 3136
rect 6125 3017 6147 3023
rect 6061 2884 6067 2916
rect 6077 2904 6083 2916
rect 6093 2864 6099 2956
rect 6045 2704 6051 2756
rect 5997 2584 6003 2616
rect 6013 2584 6019 2676
rect 5917 2557 5939 2563
rect 5885 2484 5891 2536
rect 5901 2463 5907 2556
rect 5917 2544 5923 2557
rect 6029 2544 6035 2636
rect 5933 2524 5939 2536
rect 6045 2524 6051 2676
rect 5917 2484 5923 2496
rect 5933 2464 5939 2496
rect 5892 2457 5907 2463
rect 5853 2304 5859 2356
rect 5869 2284 5875 2336
rect 5885 2324 5891 2456
rect 5901 2404 5907 2436
rect 5869 2184 5875 2276
rect 5837 2177 5859 2183
rect 5837 2124 5843 2136
rect 5853 1983 5859 2177
rect 5885 2163 5891 2236
rect 5869 2157 5891 2163
rect 5869 2104 5875 2157
rect 5885 2104 5891 2136
rect 5885 2084 5891 2096
rect 5837 1977 5859 1983
rect 5789 1784 5795 1836
rect 5629 1744 5635 1776
rect 5709 1764 5715 1776
rect 5693 1544 5699 1556
rect 5709 1544 5715 1716
rect 5725 1704 5731 1736
rect 5805 1704 5811 1856
rect 5821 1804 5827 1836
rect 5837 1783 5843 1977
rect 5853 1944 5859 1956
rect 5869 1904 5875 2076
rect 5901 2004 5907 2376
rect 5917 2304 5923 2336
rect 5949 2283 5955 2476
rect 5917 2277 5955 2283
rect 5917 1923 5923 2277
rect 5940 2257 5955 2263
rect 5933 2124 5939 2236
rect 5949 2184 5955 2257
rect 5949 2164 5955 2176
rect 5933 1964 5939 2096
rect 5965 1984 5971 2436
rect 5981 2323 5987 2496
rect 5997 2404 6003 2516
rect 6029 2497 6044 2503
rect 5997 2344 6003 2376
rect 6029 2364 6035 2497
rect 6061 2404 6067 2856
rect 6077 2524 6083 2596
rect 6093 2583 6099 2696
rect 6109 2684 6115 2916
rect 6125 2804 6131 2876
rect 6125 2704 6131 2716
rect 6141 2684 6147 3017
rect 6157 2944 6163 3056
rect 6157 2924 6163 2936
rect 6173 2824 6179 2896
rect 6157 2684 6163 2716
rect 6173 2704 6179 2716
rect 6093 2577 6115 2583
rect 6109 2564 6115 2577
rect 6093 2483 6099 2556
rect 6093 2477 6115 2483
rect 6077 2384 6083 2416
rect 5981 2317 6003 2323
rect 5981 2244 5987 2256
rect 5981 2144 5987 2216
rect 5981 1924 5987 2116
rect 5997 2023 6003 2317
rect 6013 2304 6019 2356
rect 6013 2184 6019 2276
rect 6029 2204 6035 2336
rect 6013 2144 6019 2176
rect 6029 2144 6035 2196
rect 6045 2144 6051 2316
rect 6077 2284 6083 2296
rect 6013 2043 6019 2116
rect 6029 2104 6035 2136
rect 6045 2084 6051 2116
rect 6061 2104 6067 2236
rect 6077 2204 6083 2276
rect 6093 2143 6099 2456
rect 6109 2344 6115 2477
rect 6125 2303 6131 2676
rect 6141 2424 6147 2636
rect 6157 2584 6163 2616
rect 6157 2524 6163 2576
rect 6157 2384 6163 2496
rect 6173 2304 6179 2676
rect 6189 2624 6195 2876
rect 6205 2744 6211 3056
rect 6237 2944 6243 3036
rect 6221 2784 6227 2816
rect 6237 2784 6243 2936
rect 6205 2684 6211 2696
rect 6189 2524 6195 2576
rect 6189 2364 6195 2436
rect 6109 2297 6131 2303
rect 6109 2184 6115 2297
rect 6141 2204 6147 2236
rect 6093 2137 6115 2143
rect 6013 2037 6051 2043
rect 5997 2017 6019 2023
rect 5917 1917 5955 1923
rect 5901 1864 5907 1916
rect 5917 1884 5923 1896
rect 5885 1784 5891 1856
rect 5821 1777 5843 1783
rect 5716 1537 5731 1543
rect 5725 1524 5731 1537
rect 5581 1384 5587 1396
rect 5629 1324 5635 1336
rect 5645 1323 5651 1456
rect 5709 1444 5715 1516
rect 5725 1504 5731 1516
rect 5741 1504 5747 1616
rect 5821 1524 5827 1777
rect 5917 1744 5923 1816
rect 5933 1804 5939 1896
rect 5949 1764 5955 1917
rect 5965 1844 5971 1916
rect 5981 1884 5987 1896
rect 5837 1544 5843 1676
rect 5853 1664 5859 1716
rect 5837 1524 5843 1536
rect 5853 1504 5859 1656
rect 5949 1584 5955 1716
rect 5981 1704 5987 1718
rect 5741 1484 5747 1496
rect 5821 1484 5827 1496
rect 5773 1444 5779 1456
rect 5661 1324 5667 1356
rect 5773 1324 5779 1436
rect 5645 1317 5660 1323
rect 5613 1284 5619 1316
rect 5645 1304 5651 1317
rect 5181 1164 5187 1236
rect 5133 1064 5139 1116
rect 4909 984 4915 1036
rect 4589 964 4595 976
rect 4605 957 4620 963
rect 4157 937 4179 943
rect 4157 924 4163 937
rect 4605 943 4611 957
rect 4749 944 4755 956
rect 4877 944 4883 976
rect 4596 937 4611 943
rect 4125 697 4147 703
rect 4125 684 4131 697
rect 4173 684 4179 916
rect 4237 904 4243 936
rect 4573 924 4579 936
rect 4461 904 4467 916
rect 4925 904 4931 936
rect 4957 924 4963 936
rect 3917 564 3923 636
rect 3949 543 3955 596
rect 3940 537 3955 543
rect 3869 524 3875 536
rect 3853 517 3868 523
rect 3853 464 3859 517
rect 3869 484 3875 496
rect 3901 484 3907 536
rect 3965 524 3971 536
rect 3949 484 3955 496
rect 3981 484 3987 556
rect 4013 544 4019 676
rect 4189 644 4195 656
rect 4013 504 4019 536
rect 4029 483 4035 516
rect 4045 484 4051 576
rect 4013 477 4035 483
rect 3389 284 3395 296
rect 3501 264 3507 296
rect 3533 264 3539 336
rect 3661 324 3667 336
rect 3533 243 3539 256
rect 3517 237 3539 243
rect 3112 206 3118 214
rect 3126 206 3132 214
rect 3140 206 3146 214
rect 3154 206 3160 214
rect 3517 184 3523 237
rect 3597 204 3603 296
rect 2724 157 2739 163
rect 2605 144 2611 156
rect 2733 143 2739 157
rect 2813 144 2819 156
rect 2733 137 2787 143
rect 2509 -23 2515 16
rect 2589 -23 2595 136
rect 2653 104 2659 136
rect 2701 124 2707 136
rect 2781 104 2787 137
rect 2781 -23 2787 56
rect 2845 -23 2851 156
rect 2893 124 2899 156
rect 2893 -23 2899 116
rect 2957 -17 2963 156
rect 2973 104 2979 116
rect 2941 -23 2963 -17
rect 3021 -17 3027 136
rect 3069 104 3075 116
rect 3181 104 3187 116
rect 3053 -17 3059 96
rect 3021 -23 3043 -17
rect 3053 -23 3075 -17
rect 3229 -23 3235 136
rect 3261 -23 3267 96
rect 3373 -23 3379 -17
rect 3437 -23 3443 56
rect 3485 -17 3491 156
rect 3501 144 3507 156
rect 3501 24 3507 136
rect 3533 104 3539 196
rect 3613 184 3619 196
rect 3645 164 3651 256
rect 3677 184 3683 416
rect 3693 384 3699 396
rect 3885 384 3891 456
rect 4013 404 4019 477
rect 4029 404 4035 436
rect 3789 304 3795 356
rect 3837 324 3843 356
rect 3805 264 3811 276
rect 3901 264 3907 396
rect 3933 344 3939 376
rect 3949 344 3955 356
rect 3981 304 3987 376
rect 4029 324 4035 396
rect 4045 324 4051 356
rect 3949 284 3955 296
rect 3997 284 4003 316
rect 4093 304 4099 636
rect 4109 504 4115 576
rect 4125 524 4131 536
rect 4157 464 4163 536
rect 4173 443 4179 576
rect 4189 524 4195 536
rect 4205 524 4211 656
rect 4237 584 4243 896
rect 4461 784 4467 896
rect 4372 717 4387 723
rect 4253 704 4259 716
rect 4269 584 4275 676
rect 4285 584 4291 716
rect 4301 664 4307 716
rect 4157 437 4179 443
rect 4141 384 4147 436
rect 3741 143 3747 256
rect 3773 224 3779 236
rect 3901 204 3907 256
rect 4109 204 4115 316
rect 4141 304 4147 316
rect 4141 244 4147 276
rect 4013 184 4019 196
rect 4157 184 4163 437
rect 4221 424 4227 496
rect 4237 404 4243 536
rect 4253 424 4259 516
rect 4285 384 4291 556
rect 4317 524 4323 636
rect 4333 564 4339 676
rect 4381 664 4387 717
rect 4557 704 4563 736
rect 4445 684 4451 696
rect 4381 644 4387 656
rect 4397 584 4403 636
rect 4477 584 4483 696
rect 4301 504 4307 516
rect 4381 444 4387 536
rect 4461 524 4467 556
rect 4429 444 4435 496
rect 4461 484 4467 516
rect 4493 504 4499 676
rect 4365 384 4371 416
rect 4349 324 4355 336
rect 4365 304 4371 336
rect 4276 297 4291 303
rect 4253 244 4259 276
rect 4285 263 4291 297
rect 4429 284 4435 316
rect 4461 304 4467 436
rect 4525 424 4531 696
rect 4541 684 4547 696
rect 4573 684 4579 716
rect 4605 704 4611 836
rect 4632 806 4638 814
rect 4646 806 4652 814
rect 4660 806 4666 814
rect 4674 806 4680 814
rect 4845 784 4851 896
rect 4925 884 4931 896
rect 4813 724 4819 756
rect 4845 724 4851 776
rect 4973 764 4979 1036
rect 4989 984 4995 1036
rect 5037 984 5043 996
rect 5053 964 5059 976
rect 5021 944 5027 956
rect 5053 784 5059 936
rect 5069 924 5075 1036
rect 5117 984 5123 1036
rect 5085 884 5091 976
rect 5101 904 5107 916
rect 5117 904 5123 956
rect 5133 944 5139 1016
rect 5149 964 5155 1056
rect 5197 1044 5203 1096
rect 5261 1064 5267 1136
rect 5325 1084 5331 1236
rect 5341 1124 5347 1136
rect 5245 1024 5251 1036
rect 5277 984 5283 1056
rect 5293 1044 5299 1076
rect 5341 1063 5347 1116
rect 5373 1104 5379 1136
rect 5332 1057 5347 1063
rect 5357 1044 5363 1096
rect 5405 1044 5411 1056
rect 5293 984 5299 1036
rect 5309 984 5315 1036
rect 5437 1004 5443 1076
rect 5485 1024 5491 1116
rect 5581 1084 5587 1096
rect 5517 1064 5523 1076
rect 5661 1064 5667 1096
rect 5485 984 5491 996
rect 5149 924 5155 936
rect 5101 864 5107 876
rect 5165 724 5171 916
rect 5181 904 5187 976
rect 5405 944 5411 976
rect 5181 884 5187 896
rect 5197 844 5203 936
rect 5341 924 5347 936
rect 5501 924 5507 1036
rect 5229 904 5235 916
rect 5469 864 5475 916
rect 5341 744 5347 756
rect 5293 724 5299 736
rect 4909 704 4915 716
rect 4916 697 4931 703
rect 4541 624 4547 656
rect 4557 504 4563 576
rect 4573 424 4579 676
rect 4605 664 4611 696
rect 4829 664 4835 696
rect 4877 664 4883 696
rect 4925 664 4931 697
rect 4957 664 4963 676
rect 4717 564 4723 616
rect 4589 504 4595 536
rect 4717 504 4723 556
rect 4765 544 4771 576
rect 4749 504 4755 516
rect 4765 484 4771 536
rect 4797 524 4803 616
rect 4845 577 4876 583
rect 4845 564 4851 577
rect 4861 504 4867 556
rect 4541 384 4547 416
rect 4632 406 4638 414
rect 4646 406 4652 414
rect 4660 406 4666 414
rect 4674 406 4680 414
rect 4909 344 4915 636
rect 4957 564 4963 596
rect 4973 584 4979 616
rect 4973 504 4979 536
rect 5021 484 5027 716
rect 5053 644 5059 696
rect 5085 684 5091 716
rect 5069 664 5075 676
rect 5117 644 5123 716
rect 5437 704 5443 716
rect 5453 704 5459 836
rect 5517 804 5523 936
rect 5533 904 5539 1056
rect 5549 984 5555 1016
rect 5581 964 5587 1036
rect 5629 1024 5635 1056
rect 5645 964 5651 1036
rect 5677 1024 5683 1056
rect 5581 924 5587 956
rect 5645 904 5651 956
rect 5677 924 5683 936
rect 5549 864 5555 896
rect 5629 864 5635 896
rect 5661 884 5667 916
rect 5565 744 5571 836
rect 5069 363 5075 456
rect 5085 444 5091 556
rect 5117 544 5123 576
rect 5133 524 5139 536
rect 5165 524 5171 576
rect 5181 523 5187 636
rect 5197 624 5203 696
rect 5213 684 5219 696
rect 5341 684 5347 696
rect 5213 624 5219 676
rect 5373 664 5379 696
rect 5469 684 5475 736
rect 5533 724 5539 736
rect 5517 704 5523 716
rect 5501 684 5507 696
rect 5549 684 5555 696
rect 5197 544 5203 616
rect 5213 564 5219 576
rect 5181 517 5203 523
rect 5101 464 5107 516
rect 5133 504 5139 516
rect 5149 444 5155 496
rect 5181 484 5187 496
rect 5101 384 5107 416
rect 5069 357 5091 363
rect 4477 324 4483 336
rect 4484 317 4499 323
rect 4445 264 4451 296
rect 4493 264 4499 317
rect 4781 304 4787 316
rect 4877 284 4883 296
rect 4525 264 4531 276
rect 4276 257 4291 263
rect 4260 237 4275 243
rect 3725 137 3747 143
rect 3549 124 3555 136
rect 3661 104 3667 116
rect 3709 104 3715 116
rect 3533 44 3539 96
rect 3469 -23 3491 -17
rect 3533 -23 3539 16
rect 3565 -23 3571 36
rect 3725 -23 3731 137
rect 3757 -17 3763 136
rect 3933 124 3939 156
rect 3796 97 3811 103
rect 3757 -23 3779 -17
rect 3805 -23 3811 97
rect 4077 -17 4083 156
rect 4061 -23 4083 -17
rect 4125 -23 4131 36
rect 4205 -23 4211 156
rect 4269 144 4275 237
rect 4301 144 4307 156
rect 4381 144 4387 156
rect 4253 124 4259 136
rect 4253 -23 4259 36
rect 4381 -17 4387 136
rect 4429 104 4435 156
rect 4477 124 4483 236
rect 4589 224 4595 256
rect 4621 144 4627 176
rect 4749 164 4755 276
rect 4525 124 4531 136
rect 4813 124 4819 236
rect 4861 164 4867 196
rect 4877 184 4883 276
rect 4909 264 4915 296
rect 4893 164 4899 236
rect 4925 164 4931 176
rect 4957 164 4963 336
rect 5069 304 5075 336
rect 5085 303 5091 357
rect 5165 324 5171 436
rect 5085 297 5100 303
rect 5005 264 5011 276
rect 4989 203 4995 256
rect 4973 197 4995 203
rect 4973 144 4979 197
rect 4989 144 4995 176
rect 5021 123 5027 256
rect 5012 117 5027 123
rect 5037 104 5043 276
rect 5053 264 5059 276
rect 5101 184 5107 296
rect 5133 204 5139 316
rect 5149 304 5155 316
rect 5197 304 5203 517
rect 5245 404 5251 536
rect 5309 444 5315 556
rect 5325 444 5331 636
rect 5341 544 5347 616
rect 5405 564 5411 656
rect 5501 604 5507 636
rect 5357 524 5363 536
rect 5389 504 5395 516
rect 5405 504 5411 556
rect 5469 484 5475 536
rect 5485 524 5491 556
rect 5501 504 5507 516
rect 5517 484 5523 516
rect 5533 484 5539 556
rect 5581 544 5587 636
rect 5693 584 5699 1156
rect 5709 1004 5715 1056
rect 5709 704 5715 716
rect 5693 564 5699 576
rect 5645 524 5651 536
rect 5213 184 5219 276
rect 5229 264 5235 296
rect 5245 284 5251 356
rect 5261 344 5267 436
rect 5341 304 5347 316
rect 5357 284 5363 396
rect 5389 264 5395 316
rect 5421 304 5427 396
rect 5437 364 5443 436
rect 5565 424 5571 496
rect 5581 484 5587 516
rect 5629 504 5635 516
rect 5597 484 5603 496
rect 5501 284 5507 296
rect 5533 284 5539 296
rect 5549 284 5555 336
rect 5581 324 5587 436
rect 5613 404 5619 476
rect 5677 424 5683 556
rect 5757 544 5763 1316
rect 5805 1304 5811 1436
rect 5853 1304 5859 1356
rect 5869 1344 5875 1396
rect 5901 1384 5907 1516
rect 5933 1484 5939 1536
rect 5997 1504 6003 1776
rect 6013 1684 6019 2017
rect 6029 1924 6035 2016
rect 6029 1864 6035 1876
rect 6029 1824 6035 1836
rect 6045 1744 6051 2037
rect 6061 2004 6067 2096
rect 6077 2084 6083 2116
rect 6093 2084 6099 2096
rect 6109 2044 6115 2137
rect 6077 2004 6083 2036
rect 6061 1884 6067 1956
rect 6109 1904 6115 1976
rect 6125 1964 6131 2116
rect 6141 2024 6147 2136
rect 6157 1883 6163 2236
rect 6173 2124 6179 2216
rect 6189 2144 6195 2236
rect 6221 2164 6227 2716
rect 6237 2364 6243 2556
rect 6237 2284 6243 2336
rect 6253 2224 6259 4256
rect 6205 2144 6211 2156
rect 6228 2137 6243 2143
rect 6189 2124 6195 2136
rect 6173 2104 6179 2116
rect 6221 2063 6227 2116
rect 6205 2057 6227 2063
rect 6173 1924 6179 2016
rect 6141 1877 6163 1883
rect 6045 1644 6051 1716
rect 6093 1664 6099 1876
rect 6125 1683 6131 1716
rect 6116 1677 6131 1683
rect 5949 1484 5955 1496
rect 6077 1484 6083 1636
rect 6141 1504 6147 1877
rect 6164 1857 6179 1863
rect 6173 1744 6179 1857
rect 6189 1724 6195 1836
rect 6157 1684 6163 1696
rect 6205 1584 6211 2057
rect 6221 1984 6227 2036
rect 6237 2004 6243 2137
rect 6237 1864 6243 1876
rect 6253 1784 6259 2156
rect 6237 1704 6243 1736
rect 5949 1463 5955 1476
rect 5933 1457 5955 1463
rect 5933 1384 5939 1457
rect 5917 1364 5923 1376
rect 5949 1344 5955 1416
rect 5997 1364 6003 1376
rect 6077 1344 6083 1476
rect 5917 1102 5923 1116
rect 5853 1064 5859 1076
rect 5789 904 5795 956
rect 5917 924 5923 1056
rect 5949 943 5955 1336
rect 6013 1324 6019 1336
rect 6013 1264 6019 1296
rect 6029 984 6035 1236
rect 6077 1084 6083 1336
rect 6109 1326 6115 1436
rect 6173 984 6179 1556
rect 6221 1237 6236 1243
rect 6093 944 6099 976
rect 6157 964 6163 976
rect 5949 937 5964 943
rect 5789 684 5795 896
rect 5917 784 5923 916
rect 5885 704 5891 736
rect 5917 724 5923 776
rect 5789 544 5795 676
rect 5805 524 5811 596
rect 5853 564 5859 596
rect 5629 284 5635 356
rect 5645 324 5651 336
rect 5309 164 5315 176
rect 5060 137 5084 143
rect 5229 124 5235 156
rect 5261 144 5267 156
rect 5373 143 5379 236
rect 5373 137 5388 143
rect 5405 123 5411 216
rect 5437 184 5443 236
rect 5469 184 5475 256
rect 5485 183 5491 236
rect 5549 184 5555 196
rect 5485 177 5507 183
rect 5501 144 5507 177
rect 5396 117 5411 123
rect 5421 84 5427 96
rect 5549 84 5555 136
rect 5565 124 5571 236
rect 5645 164 5651 316
rect 5677 264 5683 296
rect 5661 124 5667 256
rect 5693 183 5699 276
rect 5709 264 5715 436
rect 5741 364 5747 516
rect 5773 484 5779 496
rect 5741 284 5747 356
rect 5821 344 5827 516
rect 5837 504 5843 536
rect 5869 384 5875 636
rect 5885 564 5891 676
rect 5965 644 5971 936
rect 6205 924 6211 1036
rect 6093 904 6099 916
rect 5981 884 5987 896
rect 6141 884 6147 896
rect 5997 664 6003 776
rect 6029 704 6035 836
rect 6205 784 6211 876
rect 6132 737 6147 743
rect 6141 704 6147 737
rect 6173 684 6179 696
rect 6189 684 6195 736
rect 6205 663 6211 696
rect 6221 664 6227 1237
rect 6237 1024 6243 1036
rect 6189 657 6211 663
rect 5933 584 5939 636
rect 5917 544 5923 556
rect 5821 304 5827 316
rect 5741 224 5747 236
rect 5684 177 5699 183
rect 5677 144 5683 176
rect 5805 164 5811 196
rect 5709 124 5715 136
rect 5565 104 5571 116
rect 5821 84 5827 296
rect 5869 204 5875 296
rect 5901 284 5907 316
rect 5885 264 5891 276
rect 5917 244 5923 296
rect 5933 183 5939 256
rect 5949 184 5955 616
rect 5997 544 6003 656
rect 5981 243 5987 536
rect 6173 524 6179 656
rect 6036 517 6051 523
rect 6045 384 6051 517
rect 6125 483 6131 516
rect 6116 477 6131 483
rect 5997 304 6003 316
rect 6013 284 6019 336
rect 6109 264 6115 276
rect 5981 237 6003 243
rect 5917 177 5939 183
rect 5917 144 5923 177
rect 5933 144 5939 156
rect 5997 144 6003 237
rect 6125 184 6131 296
rect 6157 263 6163 436
rect 6173 304 6179 496
rect 6189 343 6195 657
rect 6221 584 6227 636
rect 6253 544 6259 1596
rect 6221 504 6227 516
rect 6205 484 6211 496
rect 6237 384 6243 456
rect 6189 337 6211 343
rect 6141 257 6163 263
rect 6029 104 6035 118
rect 4381 -23 4403 -17
rect 4429 -23 4435 76
rect 5613 64 5619 76
rect 4509 -17 4515 36
rect 4557 -17 4563 36
rect 4632 6 4638 14
rect 4646 6 4652 14
rect 4660 6 4666 14
rect 4674 6 4680 14
rect 4493 -23 4515 -17
rect 4541 -23 4563 -17
rect 4685 -23 4691 -17
rect 4845 -23 4851 16
rect 5917 -23 5923 16
rect 6109 -23 6115 -17
rect 6141 -23 6147 257
rect 6157 204 6163 236
rect 6205 184 6211 337
rect 6253 284 6259 316
rect 6173 -23 6179 16
<< m3contact >>
rect 460 5796 468 5804
rect 492 5796 500 5804
rect 60 5756 68 5764
rect 124 5756 132 5764
rect 300 5756 308 5764
rect 28 5716 36 5724
rect 124 5736 132 5744
rect 156 5736 164 5744
rect 220 5736 228 5744
rect 284 5736 292 5744
rect 364 5736 372 5744
rect 396 5736 404 5744
rect 76 5716 84 5724
rect 44 5696 52 5704
rect 76 5696 84 5704
rect 140 5716 148 5724
rect 204 5716 212 5724
rect 252 5716 260 5724
rect 444 5716 452 5724
rect 188 5596 196 5604
rect 668 5776 676 5784
rect 652 5756 660 5764
rect 540 5736 548 5744
rect 588 5736 596 5744
rect 796 5736 804 5744
rect 508 5716 516 5724
rect 540 5716 548 5724
rect 572 5716 580 5724
rect 780 5716 788 5724
rect 364 5696 372 5704
rect 396 5696 404 5704
rect 492 5696 500 5704
rect 540 5696 548 5704
rect 588 5696 596 5704
rect 828 5796 836 5804
rect 812 5716 820 5724
rect 956 5756 964 5764
rect 844 5696 852 5704
rect 316 5656 324 5664
rect 236 5596 244 5604
rect 284 5596 292 5604
rect 204 5576 212 5584
rect 44 5556 52 5564
rect 604 5676 612 5684
rect 716 5556 724 5564
rect 92 5536 100 5544
rect 236 5536 244 5544
rect 348 5536 356 5544
rect 12 5476 20 5484
rect 220 5516 228 5524
rect 268 5516 276 5524
rect 188 5496 196 5504
rect 12 5376 20 5384
rect 28 5376 36 5384
rect 28 5336 36 5344
rect 44 5316 52 5324
rect 172 5476 180 5484
rect 204 5456 212 5464
rect 140 5436 148 5444
rect 172 5396 180 5404
rect 140 5356 148 5364
rect 76 5296 84 5304
rect 28 5236 36 5244
rect 60 5236 68 5244
rect 252 5456 260 5464
rect 236 5416 244 5424
rect 220 5356 228 5364
rect 156 5316 164 5324
rect 140 5176 148 5184
rect 12 5056 20 5064
rect 76 5076 84 5084
rect 92 5056 100 5064
rect 268 5436 276 5444
rect 284 5436 292 5444
rect 252 5336 260 5344
rect 284 5336 292 5344
rect 252 5296 260 5304
rect 236 5236 244 5244
rect 748 5576 756 5584
rect 732 5536 740 5544
rect 780 5556 788 5564
rect 380 5496 388 5504
rect 428 5496 436 5504
rect 332 5456 340 5464
rect 396 5476 404 5484
rect 444 5476 452 5484
rect 380 5436 388 5444
rect 412 5436 420 5444
rect 460 5436 468 5444
rect 348 5416 356 5424
rect 444 5416 452 5424
rect 348 5396 356 5404
rect 444 5376 452 5384
rect 300 5316 308 5324
rect 268 5116 276 5124
rect 220 5096 228 5104
rect 188 5036 196 5044
rect 284 5096 292 5104
rect 268 5076 276 5084
rect 428 5336 436 5344
rect 492 5496 500 5504
rect 668 5496 676 5504
rect 604 5476 612 5484
rect 716 5476 724 5484
rect 508 5456 516 5464
rect 620 5456 628 5464
rect 524 5436 532 5444
rect 588 5436 596 5444
rect 492 5356 500 5364
rect 540 5416 548 5424
rect 604 5396 612 5404
rect 796 5476 804 5484
rect 796 5456 804 5464
rect 844 5676 852 5684
rect 1068 5796 1076 5804
rect 1132 5796 1140 5804
rect 1020 5776 1028 5784
rect 1084 5776 1092 5784
rect 956 5736 964 5744
rect 1020 5736 1028 5744
rect 1052 5736 1060 5744
rect 924 5696 932 5704
rect 956 5696 964 5704
rect 972 5676 980 5684
rect 908 5636 916 5644
rect 844 5576 852 5584
rect 908 5536 916 5544
rect 1004 5716 1012 5724
rect 988 5536 996 5544
rect 876 5496 884 5504
rect 940 5496 948 5504
rect 956 5496 964 5504
rect 988 5496 996 5504
rect 1020 5636 1028 5644
rect 1148 5756 1156 5764
rect 1196 5756 1204 5764
rect 1116 5736 1124 5744
rect 1132 5736 1140 5744
rect 1132 5696 1140 5704
rect 1212 5696 1220 5704
rect 1084 5656 1092 5664
rect 1100 5656 1108 5664
rect 1068 5636 1076 5644
rect 1148 5636 1156 5644
rect 1212 5636 1220 5644
rect 1052 5596 1060 5604
rect 1020 5516 1028 5524
rect 1052 5516 1060 5524
rect 908 5456 916 5464
rect 1004 5436 1012 5444
rect 988 5416 996 5424
rect 828 5396 836 5404
rect 1004 5396 1012 5404
rect 652 5376 660 5384
rect 844 5376 852 5384
rect 1164 5596 1172 5604
rect 1100 5576 1108 5584
rect 1116 5456 1124 5464
rect 1148 5456 1156 5464
rect 1148 5436 1156 5444
rect 1100 5396 1108 5404
rect 1132 5376 1140 5384
rect 716 5356 724 5364
rect 1068 5356 1076 5364
rect 1132 5356 1140 5364
rect 492 5336 500 5344
rect 540 5336 548 5344
rect 412 5316 420 5324
rect 444 5316 452 5324
rect 396 5296 404 5304
rect 396 5236 404 5244
rect 380 5116 388 5124
rect 332 5096 340 5104
rect 316 5056 324 5064
rect 252 5036 260 5044
rect 364 5056 372 5064
rect 380 5036 388 5044
rect 556 5316 564 5324
rect 620 5316 628 5324
rect 444 5296 452 5304
rect 476 5296 484 5304
rect 508 5296 516 5304
rect 428 5096 436 5104
rect 476 5096 484 5104
rect 444 5076 452 5084
rect 444 5056 452 5064
rect 492 5076 500 5084
rect 572 5296 580 5304
rect 636 5276 644 5284
rect 732 5336 740 5344
rect 844 5336 852 5344
rect 828 5316 836 5324
rect 892 5316 900 5324
rect 828 5176 836 5184
rect 1036 5316 1044 5324
rect 1068 5316 1076 5324
rect 1116 5316 1124 5324
rect 1292 5796 1300 5804
rect 1388 5736 1396 5744
rect 1404 5736 1412 5744
rect 1324 5696 1332 5704
rect 1292 5616 1300 5624
rect 1340 5616 1348 5624
rect 3118 5806 3126 5814
rect 3132 5806 3140 5814
rect 3146 5806 3154 5814
rect 1548 5796 1556 5804
rect 3036 5796 3044 5804
rect 1468 5716 1476 5724
rect 1420 5676 1428 5684
rect 1452 5676 1460 5684
rect 1372 5656 1380 5664
rect 1356 5596 1364 5604
rect 1372 5596 1380 5604
rect 1340 5536 1348 5544
rect 1356 5536 1364 5544
rect 1228 5516 1236 5524
rect 1292 5516 1300 5524
rect 1276 5496 1284 5504
rect 1292 5476 1300 5484
rect 1276 5456 1284 5464
rect 1260 5396 1268 5404
rect 1244 5376 1252 5384
rect 1196 5356 1204 5364
rect 1212 5336 1220 5344
rect 1180 5316 1188 5324
rect 1084 5296 1092 5304
rect 1164 5296 1172 5304
rect 1052 5256 1060 5264
rect 828 5136 836 5144
rect 892 5136 900 5144
rect 588 5116 596 5124
rect 716 5116 724 5124
rect 764 5116 772 5124
rect 956 5116 964 5124
rect 1036 5116 1044 5124
rect 700 5096 708 5104
rect 748 5076 756 5084
rect 556 4976 564 4984
rect 76 4956 84 4964
rect 220 4956 228 4964
rect 108 4936 116 4944
rect 76 4796 84 4804
rect 828 5096 836 5104
rect 860 5096 868 5104
rect 956 5096 964 5104
rect 924 5076 932 5084
rect 732 5056 740 5064
rect 780 5056 788 5064
rect 892 5056 900 5064
rect 940 5056 948 5064
rect 940 5016 948 5024
rect 1004 5096 1012 5104
rect 988 5076 996 5084
rect 1004 5056 1012 5064
rect 924 4976 932 4984
rect 732 4956 740 4964
rect 956 4956 964 4964
rect 364 4936 372 4944
rect 412 4936 420 4944
rect 492 4936 500 4944
rect 524 4936 532 4944
rect 844 4936 852 4944
rect 988 4936 996 4944
rect 156 4916 164 4924
rect 204 4916 212 4924
rect 316 4916 324 4924
rect 124 4896 132 4904
rect 172 4896 180 4904
rect 124 4796 132 4804
rect 188 4696 196 4704
rect 156 4680 164 4684
rect 156 4676 164 4680
rect 12 4656 20 4664
rect 76 4636 84 4644
rect 108 4596 116 4604
rect 124 4556 132 4564
rect 76 4516 84 4524
rect 12 4456 20 4464
rect 44 4376 52 4384
rect 12 4336 20 4344
rect 60 4296 68 4304
rect 44 4276 52 4284
rect 188 4556 196 4564
rect 284 4896 292 4904
rect 332 4896 340 4904
rect 380 4896 388 4904
rect 668 4916 676 4924
rect 508 4896 516 4904
rect 556 4896 564 4904
rect 700 4896 708 4904
rect 764 4916 772 4924
rect 892 4916 900 4924
rect 940 4896 948 4904
rect 748 4856 756 4864
rect 716 4816 724 4824
rect 780 4816 788 4824
rect 636 4716 644 4724
rect 684 4716 692 4724
rect 332 4696 340 4704
rect 476 4696 484 4704
rect 236 4676 244 4684
rect 444 4676 452 4684
rect 220 4596 228 4604
rect 108 4436 116 4444
rect 172 4316 180 4324
rect 92 4276 100 4284
rect 108 4276 116 4284
rect 140 4276 148 4284
rect 236 4536 244 4544
rect 236 4396 244 4404
rect 204 4336 212 4344
rect 220 4316 228 4324
rect 220 4296 228 4304
rect 268 4636 276 4644
rect 444 4656 452 4664
rect 476 4656 484 4664
rect 268 4616 276 4624
rect 348 4616 356 4624
rect 508 4656 516 4664
rect 668 4696 676 4704
rect 940 4736 948 4744
rect 892 4716 900 4724
rect 972 4716 980 4724
rect 940 4696 948 4704
rect 972 4696 980 4704
rect 844 4676 852 4684
rect 556 4656 564 4664
rect 668 4656 676 4664
rect 492 4636 500 4644
rect 524 4636 532 4644
rect 652 4636 660 4644
rect 620 4616 628 4624
rect 348 4576 356 4584
rect 492 4576 500 4584
rect 460 4536 468 4544
rect 284 4516 292 4524
rect 284 4456 292 4464
rect 268 4376 276 4384
rect 268 4236 276 4244
rect 380 4336 388 4344
rect 412 4516 420 4524
rect 476 4516 484 4524
rect 444 4496 452 4504
rect 476 4496 484 4504
rect 460 4476 468 4484
rect 572 4556 580 4564
rect 636 4556 644 4564
rect 556 4496 564 4504
rect 604 4496 612 4504
rect 540 4476 548 4484
rect 588 4476 596 4484
rect 556 4456 564 4464
rect 572 4356 580 4364
rect 412 4336 420 4344
rect 316 4296 324 4304
rect 348 4276 356 4284
rect 108 4136 116 4144
rect 220 4136 228 4144
rect 12 4116 20 4124
rect 124 4116 132 4124
rect 76 4016 84 4024
rect 124 3936 132 3944
rect 108 3896 116 3904
rect 12 3836 20 3844
rect 44 3836 52 3844
rect 188 4056 196 4064
rect 204 3936 212 3944
rect 124 3816 132 3824
rect 76 3716 84 3724
rect 12 3696 20 3704
rect 140 3736 148 3744
rect 124 3696 132 3704
rect 140 3536 148 3544
rect 172 3876 180 3884
rect 172 3816 180 3824
rect 268 4116 276 4124
rect 236 4096 244 4104
rect 236 4076 244 4084
rect 284 4056 292 4064
rect 268 3916 276 3924
rect 236 3896 244 3904
rect 252 3876 260 3884
rect 252 3856 260 3864
rect 236 3836 244 3844
rect 220 3796 228 3804
rect 188 3736 196 3744
rect 236 3716 244 3724
rect 172 3696 180 3704
rect 220 3696 228 3704
rect 188 3596 196 3604
rect 156 3496 164 3504
rect 172 3496 180 3504
rect 12 3436 20 3444
rect 44 3296 52 3304
rect 44 3256 52 3264
rect 124 3376 132 3384
rect 172 3356 180 3364
rect 300 3736 308 3744
rect 364 4256 372 4264
rect 428 4316 436 4324
rect 476 4336 484 4344
rect 572 4336 580 4344
rect 460 4296 468 4304
rect 444 4276 452 4284
rect 508 4276 516 4284
rect 652 4476 660 4484
rect 604 4336 612 4344
rect 604 4296 612 4304
rect 460 4236 468 4244
rect 492 4196 500 4204
rect 540 4156 548 4164
rect 332 4136 340 4144
rect 396 4136 404 4144
rect 332 4016 340 4024
rect 332 3996 340 4004
rect 380 4096 388 4104
rect 444 4056 452 4064
rect 428 4036 436 4044
rect 364 3936 372 3944
rect 412 3916 420 3924
rect 364 3896 372 3904
rect 396 3896 404 3904
rect 348 3856 356 3864
rect 412 3836 420 3844
rect 412 3816 420 3824
rect 380 3796 388 3804
rect 396 3756 404 3764
rect 316 3716 324 3724
rect 332 3696 340 3704
rect 300 3636 308 3644
rect 268 3596 276 3604
rect 284 3596 292 3604
rect 332 3596 340 3604
rect 268 3536 276 3544
rect 252 3516 260 3524
rect 156 3336 164 3344
rect 220 3336 228 3344
rect 124 3216 132 3224
rect 172 3216 180 3224
rect 204 3216 212 3224
rect 220 3196 228 3204
rect 412 3696 420 3704
rect 364 3656 372 3664
rect 412 3656 420 3664
rect 364 3616 372 3624
rect 396 3596 404 3604
rect 348 3576 356 3584
rect 364 3556 372 3564
rect 268 3476 276 3484
rect 348 3416 356 3424
rect 380 3496 388 3504
rect 492 4016 500 4024
rect 588 4276 596 4284
rect 636 4256 644 4264
rect 588 4216 596 4224
rect 604 4156 612 4164
rect 652 4156 660 4164
rect 588 4136 596 4144
rect 620 4096 628 4104
rect 588 4036 596 4044
rect 588 3956 596 3964
rect 556 3936 564 3944
rect 476 3896 484 3904
rect 444 3816 452 3824
rect 460 3756 468 3764
rect 476 3736 484 3744
rect 476 3716 484 3724
rect 460 3696 468 3704
rect 476 3656 484 3664
rect 444 3636 452 3644
rect 428 3616 436 3624
rect 476 3596 484 3604
rect 780 4636 788 4644
rect 876 4616 884 4624
rect 828 4596 836 4604
rect 892 4596 900 4604
rect 860 4576 868 4584
rect 972 4576 980 4584
rect 1068 5136 1076 5144
rect 1100 5096 1108 5104
rect 1068 5076 1076 5084
rect 1052 5056 1060 5064
rect 1052 5036 1060 5044
rect 1100 5036 1108 5044
rect 1084 4996 1092 5004
rect 1068 4956 1076 4964
rect 1036 4916 1044 4924
rect 1100 4936 1108 4944
rect 1020 4896 1028 4904
rect 1068 4896 1076 4904
rect 1084 4896 1092 4904
rect 1036 4876 1044 4884
rect 1196 5296 1204 5304
rect 1180 5136 1188 5144
rect 1244 5116 1252 5124
rect 1180 5056 1188 5064
rect 1164 5036 1172 5044
rect 1132 5016 1140 5024
rect 1164 4996 1172 5004
rect 1420 5576 1428 5584
rect 1436 5536 1444 5544
rect 3228 5776 3236 5784
rect 3356 5776 3364 5784
rect 3420 5776 3428 5784
rect 1596 5756 1604 5764
rect 1772 5756 1780 5764
rect 1820 5756 1828 5764
rect 1852 5756 1860 5764
rect 1932 5756 1940 5764
rect 1964 5756 1972 5764
rect 1980 5756 1988 5764
rect 2156 5756 2164 5764
rect 2220 5756 2228 5764
rect 2668 5756 2676 5764
rect 2716 5756 2724 5764
rect 2780 5756 2788 5764
rect 3020 5756 3028 5764
rect 1628 5716 1636 5724
rect 1644 5716 1652 5724
rect 1516 5696 1524 5704
rect 1500 5596 1508 5604
rect 1566 5606 1574 5614
rect 1580 5606 1588 5614
rect 1594 5606 1602 5614
rect 1516 5576 1524 5584
rect 1548 5576 1556 5584
rect 1580 5576 1588 5584
rect 1452 5516 1460 5524
rect 1468 5516 1476 5524
rect 1388 5496 1396 5504
rect 1404 5496 1412 5504
rect 1340 5456 1348 5464
rect 1388 5456 1396 5464
rect 1324 5436 1332 5444
rect 1308 5336 1316 5344
rect 1420 5336 1428 5344
rect 1308 5316 1316 5324
rect 1356 5316 1364 5324
rect 1420 5316 1428 5324
rect 1340 5296 1348 5304
rect 1292 5276 1300 5284
rect 1324 5116 1332 5124
rect 1372 5276 1380 5284
rect 1404 5276 1412 5284
rect 1580 5496 1588 5504
rect 1612 5496 1620 5504
rect 1484 5476 1492 5484
rect 1468 5416 1476 5424
rect 1468 5316 1476 5324
rect 1452 5296 1460 5304
rect 1484 5296 1492 5304
rect 1516 5476 1524 5484
rect 1532 5436 1540 5444
rect 1724 5736 1732 5744
rect 1676 5696 1684 5704
rect 1708 5676 1716 5684
rect 1756 5676 1764 5684
rect 1772 5656 1780 5664
rect 1804 5676 1812 5684
rect 1900 5736 1908 5744
rect 2092 5736 2100 5744
rect 2124 5736 2132 5744
rect 1916 5716 1924 5724
rect 1932 5716 1940 5724
rect 1996 5716 2004 5724
rect 1868 5696 1876 5704
rect 2028 5716 2036 5724
rect 2044 5716 2052 5724
rect 2140 5716 2148 5724
rect 2204 5716 2212 5724
rect 2300 5716 2308 5724
rect 2332 5716 2340 5724
rect 2076 5696 2084 5704
rect 2188 5696 2196 5704
rect 2252 5696 2260 5704
rect 1884 5676 1892 5684
rect 1948 5676 1956 5684
rect 2044 5676 2052 5684
rect 2060 5676 2068 5684
rect 2124 5676 2132 5684
rect 2268 5676 2276 5684
rect 2652 5736 2660 5744
rect 2700 5736 2708 5744
rect 2796 5736 2804 5744
rect 3212 5736 3220 5744
rect 2348 5696 2356 5704
rect 2364 5696 2372 5704
rect 2396 5676 2404 5684
rect 2412 5676 2420 5684
rect 2284 5656 2292 5664
rect 2380 5656 2388 5664
rect 1788 5616 1796 5624
rect 1852 5616 1860 5624
rect 1916 5616 1924 5624
rect 1884 5576 1892 5584
rect 2204 5576 2212 5584
rect 1980 5536 1988 5544
rect 2044 5536 2052 5544
rect 2140 5536 2148 5544
rect 1932 5516 1940 5524
rect 1772 5496 1780 5504
rect 1660 5476 1668 5484
rect 1692 5476 1700 5484
rect 1628 5456 1636 5464
rect 1708 5436 1716 5444
rect 1628 5416 1636 5424
rect 1644 5416 1652 5424
rect 1612 5356 1620 5364
rect 1532 5336 1540 5344
rect 1500 5276 1508 5284
rect 1516 5276 1524 5284
rect 1596 5296 1604 5304
rect 1436 5256 1444 5264
rect 1564 5256 1572 5264
rect 1436 5236 1444 5244
rect 1372 5096 1380 5104
rect 1420 5096 1428 5104
rect 1292 5076 1300 5084
rect 1212 4996 1220 5004
rect 1196 4956 1204 4964
rect 1148 4936 1156 4944
rect 1148 4916 1156 4924
rect 1244 5016 1252 5024
rect 1356 5056 1364 5064
rect 1308 5036 1316 5044
rect 1420 5056 1428 5064
rect 1420 5016 1428 5024
rect 1244 4996 1252 5004
rect 1276 4996 1284 5004
rect 1372 4996 1380 5004
rect 1228 4976 1236 4984
rect 1212 4916 1220 4924
rect 1164 4876 1172 4884
rect 1116 4796 1124 4804
rect 1052 4696 1060 4704
rect 1084 4676 1092 4684
rect 1164 4676 1172 4684
rect 1020 4656 1028 4664
rect 1132 4656 1140 4664
rect 1164 4656 1172 4664
rect 1180 4656 1188 4664
rect 988 4556 996 4564
rect 1020 4636 1028 4644
rect 1100 4596 1108 4604
rect 1244 4956 1252 4964
rect 1372 4956 1380 4964
rect 1566 5206 1574 5214
rect 1580 5206 1588 5214
rect 1594 5206 1602 5214
rect 1468 5116 1476 5124
rect 1644 5336 1652 5344
rect 2108 5516 2116 5524
rect 1756 5476 1764 5484
rect 2092 5476 2100 5484
rect 1788 5436 1796 5444
rect 1836 5436 1844 5444
rect 1692 5356 1700 5364
rect 1692 5336 1700 5344
rect 1692 5316 1700 5324
rect 1724 5356 1732 5364
rect 1708 5256 1716 5264
rect 1740 5276 1748 5284
rect 1772 5276 1780 5284
rect 1756 5256 1764 5264
rect 1692 5216 1700 5224
rect 1724 5216 1732 5224
rect 1740 5116 1748 5124
rect 1772 5136 1780 5144
rect 1628 5096 1636 5104
rect 1676 5096 1684 5104
rect 1580 5076 1588 5084
rect 1724 5076 1732 5084
rect 1644 5056 1652 5064
rect 1724 5056 1732 5064
rect 1708 5036 1716 5044
rect 1596 5016 1604 5024
rect 1260 4936 1268 4944
rect 1356 4936 1364 4944
rect 1404 4936 1412 4944
rect 1324 4916 1332 4924
rect 1308 4876 1316 4884
rect 1372 4816 1380 4824
rect 1324 4796 1332 4804
rect 1404 4776 1412 4784
rect 1292 4756 1300 4764
rect 1324 4736 1332 4744
rect 1388 4736 1396 4744
rect 1276 4676 1284 4684
rect 1452 4816 1460 4824
rect 1452 4736 1460 4744
rect 1436 4716 1444 4724
rect 1308 4696 1316 4704
rect 1372 4696 1380 4704
rect 1420 4696 1428 4704
rect 1196 4636 1204 4644
rect 1228 4636 1236 4644
rect 1164 4616 1172 4624
rect 1292 4616 1300 4624
rect 1452 4676 1460 4684
rect 1516 4936 1524 4944
rect 1820 5316 1828 5324
rect 2188 5516 2196 5524
rect 2284 5576 2292 5584
rect 2364 5576 2372 5584
rect 2332 5536 2340 5544
rect 2380 5536 2388 5544
rect 2300 5516 2308 5524
rect 2172 5496 2180 5504
rect 2284 5496 2292 5504
rect 1916 5456 1924 5464
rect 1948 5456 1956 5464
rect 2092 5456 2100 5464
rect 2124 5456 2132 5464
rect 2220 5456 2228 5464
rect 1900 5436 1908 5444
rect 1868 5416 1876 5424
rect 1996 5436 2004 5444
rect 2092 5396 2100 5404
rect 2492 5696 2500 5704
rect 2428 5636 2436 5644
rect 2572 5716 2580 5724
rect 2620 5716 2628 5724
rect 2780 5716 2788 5724
rect 2684 5696 2692 5704
rect 2748 5696 2756 5704
rect 2556 5636 2564 5644
rect 2572 5636 2580 5644
rect 2540 5616 2548 5624
rect 2444 5576 2452 5584
rect 2428 5516 2436 5524
rect 2364 5496 2372 5504
rect 2396 5496 2404 5504
rect 2348 5476 2356 5484
rect 2316 5376 2324 5384
rect 2380 5456 2388 5464
rect 2428 5436 2436 5444
rect 2268 5356 2276 5364
rect 2364 5356 2372 5364
rect 2412 5356 2420 5364
rect 1868 5316 1876 5324
rect 1916 5316 1924 5324
rect 1820 5296 1828 5304
rect 1804 5276 1812 5284
rect 1900 5296 1908 5304
rect 1948 5296 1956 5304
rect 1852 5276 1860 5284
rect 1820 5096 1828 5104
rect 1820 5076 1828 5084
rect 1788 4996 1796 5004
rect 1868 5076 1876 5084
rect 1836 5056 1844 5064
rect 1852 5056 1860 5064
rect 1868 4976 1876 4984
rect 1836 4956 1844 4964
rect 2044 5336 2052 5344
rect 1980 5296 1988 5304
rect 2028 5276 2036 5284
rect 2076 5276 2084 5284
rect 2012 5256 2020 5264
rect 1964 5236 1972 5244
rect 1996 5236 2004 5244
rect 2108 5296 2116 5304
rect 2092 5256 2100 5264
rect 2140 5316 2148 5324
rect 2204 5316 2212 5324
rect 2172 5296 2180 5304
rect 2156 5276 2164 5284
rect 2188 5276 2196 5284
rect 2172 5256 2180 5264
rect 1996 5176 2004 5184
rect 1916 5116 1924 5124
rect 1916 5096 1924 5104
rect 1916 4996 1924 5004
rect 2140 5136 2148 5144
rect 1948 5116 1956 5124
rect 2332 5336 2340 5344
rect 2396 5336 2404 5344
rect 2268 5316 2276 5324
rect 2364 5316 2372 5324
rect 2316 5296 2324 5304
rect 2380 5296 2388 5304
rect 2508 5416 2516 5424
rect 2572 5616 2580 5624
rect 2620 5656 2628 5664
rect 2812 5656 2820 5664
rect 2716 5636 2724 5644
rect 2860 5636 2868 5644
rect 2636 5496 2644 5504
rect 2572 5476 2580 5484
rect 2620 5476 2628 5484
rect 2668 5476 2676 5484
rect 3084 5716 3092 5724
rect 2988 5696 2996 5704
rect 3292 5736 3300 5744
rect 3260 5716 3268 5724
rect 3548 5756 3556 5764
rect 3628 5756 3636 5764
rect 3852 5756 3860 5764
rect 4124 5756 4132 5764
rect 4172 5756 4180 5764
rect 3612 5736 3620 5744
rect 3804 5736 3812 5744
rect 3388 5716 3396 5724
rect 3516 5716 3524 5724
rect 3596 5716 3604 5724
rect 3692 5716 3700 5724
rect 3212 5696 3220 5704
rect 3292 5696 3300 5704
rect 3340 5696 3348 5704
rect 3468 5696 3476 5704
rect 3548 5696 3556 5704
rect 2924 5676 2932 5684
rect 3132 5676 3140 5684
rect 3244 5676 3252 5684
rect 3404 5676 3412 5684
rect 2748 5616 2756 5624
rect 2876 5616 2884 5624
rect 2716 5516 2724 5524
rect 3244 5556 3252 5564
rect 2860 5536 2868 5544
rect 2876 5536 2884 5544
rect 2908 5536 2916 5544
rect 2972 5536 2980 5544
rect 3004 5536 3012 5544
rect 3228 5536 3236 5544
rect 3260 5536 3268 5544
rect 2988 5516 2996 5524
rect 2588 5456 2596 5464
rect 2476 5376 2484 5384
rect 2540 5376 2548 5384
rect 2572 5376 2580 5384
rect 2684 5416 2692 5424
rect 2620 5356 2628 5364
rect 2508 5336 2516 5344
rect 2556 5316 2564 5324
rect 2748 5396 2756 5404
rect 2716 5356 2724 5364
rect 2828 5476 2836 5484
rect 2812 5456 2820 5464
rect 3116 5516 3124 5524
rect 3212 5516 3220 5524
rect 3180 5496 3188 5504
rect 2940 5476 2948 5484
rect 2860 5436 2868 5444
rect 2876 5416 2884 5424
rect 2812 5376 2820 5384
rect 2828 5376 2836 5384
rect 2796 5356 2804 5364
rect 2844 5356 2852 5364
rect 2764 5316 2772 5324
rect 2892 5356 2900 5364
rect 3276 5516 3284 5524
rect 3292 5496 3300 5504
rect 3340 5536 3348 5544
rect 3436 5536 3444 5544
rect 3356 5496 3364 5504
rect 3404 5496 3412 5504
rect 3052 5476 3060 5484
rect 3276 5476 3284 5484
rect 3308 5476 3316 5484
rect 3324 5476 3332 5484
rect 2956 5436 2964 5444
rect 3020 5436 3028 5444
rect 2924 5416 2932 5424
rect 2956 5356 2964 5364
rect 2652 5296 2660 5304
rect 2700 5296 2708 5304
rect 2780 5296 2788 5304
rect 2796 5296 2804 5304
rect 2860 5296 2868 5304
rect 2908 5296 2916 5304
rect 2940 5296 2948 5304
rect 3388 5476 3396 5484
rect 3484 5516 3492 5524
rect 3452 5496 3460 5504
rect 3436 5476 3444 5484
rect 3180 5456 3188 5464
rect 3420 5456 3428 5464
rect 3068 5416 3076 5424
rect 3118 5406 3126 5414
rect 3132 5406 3140 5414
rect 3146 5406 3154 5414
rect 3180 5376 3188 5384
rect 3100 5356 3108 5364
rect 3212 5376 3220 5384
rect 3020 5336 3028 5344
rect 3100 5336 3108 5344
rect 3196 5336 3204 5344
rect 3372 5376 3380 5384
rect 3340 5356 3348 5364
rect 3228 5336 3236 5344
rect 3260 5336 3268 5344
rect 3324 5336 3332 5344
rect 3004 5316 3012 5324
rect 3068 5316 3076 5324
rect 2284 5276 2292 5284
rect 2492 5276 2500 5284
rect 2668 5276 2676 5284
rect 2716 5276 2724 5284
rect 2764 5276 2772 5284
rect 2908 5276 2916 5284
rect 2972 5276 2980 5284
rect 2236 5236 2244 5244
rect 2252 5236 2260 5244
rect 2284 5236 2292 5244
rect 1964 5096 1972 5104
rect 1996 5096 2004 5104
rect 2060 5096 2068 5104
rect 2204 5096 2212 5104
rect 2364 5096 2372 5104
rect 2444 5096 2452 5104
rect 2060 5076 2068 5084
rect 2188 5076 2196 5084
rect 2236 5076 2244 5084
rect 2268 5076 2276 5084
rect 2044 5056 2052 5064
rect 2092 5056 2100 5064
rect 2172 5056 2180 5064
rect 1932 4976 1940 4984
rect 1900 4956 1908 4964
rect 1980 4956 1988 4964
rect 1884 4936 1892 4944
rect 1500 4896 1508 4904
rect 1548 4896 1556 4904
rect 1484 4876 1492 4884
rect 1484 4796 1492 4804
rect 1628 4876 1636 4884
rect 1566 4806 1574 4814
rect 1580 4806 1588 4814
rect 1594 4806 1602 4814
rect 1532 4756 1540 4764
rect 1612 4756 1620 4764
rect 1484 4696 1492 4704
rect 1516 4716 1524 4724
rect 1532 4676 1540 4684
rect 1468 4616 1476 4624
rect 1516 4616 1524 4624
rect 1340 4596 1348 4604
rect 1404 4596 1412 4604
rect 1436 4596 1444 4604
rect 1500 4596 1508 4604
rect 1820 4916 1828 4924
rect 1852 4916 1860 4924
rect 1724 4836 1732 4844
rect 1788 4756 1796 4764
rect 1660 4736 1668 4744
rect 1756 4736 1764 4744
rect 1772 4736 1780 4744
rect 1644 4696 1652 4704
rect 1676 4656 1684 4664
rect 1772 4656 1780 4664
rect 1628 4636 1636 4644
rect 1660 4636 1668 4644
rect 1644 4616 1652 4624
rect 1036 4576 1044 4584
rect 1324 4576 1332 4584
rect 1596 4576 1604 4584
rect 1724 4576 1732 4584
rect 1740 4576 1748 4584
rect 1100 4556 1108 4564
rect 1164 4556 1172 4564
rect 1228 4556 1236 4564
rect 1260 4556 1268 4564
rect 1324 4556 1332 4564
rect 748 4536 756 4544
rect 764 4536 772 4544
rect 876 4536 884 4544
rect 716 4516 724 4524
rect 684 4496 692 4504
rect 700 4496 708 4504
rect 764 4496 772 4504
rect 940 4496 948 4504
rect 700 4476 708 4484
rect 684 4436 692 4444
rect 684 4356 692 4364
rect 700 4316 708 4324
rect 748 4316 756 4324
rect 716 4296 724 4304
rect 732 4296 740 4304
rect 748 4256 756 4264
rect 988 4476 996 4484
rect 1036 4496 1044 4504
rect 1052 4496 1060 4504
rect 1084 4476 1092 4484
rect 1004 4456 1012 4464
rect 1068 4456 1076 4464
rect 908 4436 916 4444
rect 828 4396 836 4404
rect 844 4396 852 4404
rect 812 4316 820 4324
rect 796 4296 804 4304
rect 780 4276 788 4284
rect 780 4256 788 4264
rect 828 4256 836 4264
rect 764 4236 772 4244
rect 812 4236 820 4244
rect 684 4176 692 4184
rect 732 4176 740 4184
rect 684 4156 692 4164
rect 796 4156 804 4164
rect 732 4136 740 4144
rect 812 4116 820 4124
rect 1004 4376 1012 4384
rect 988 4356 996 4364
rect 940 4276 948 4284
rect 956 4276 964 4284
rect 844 4236 852 4244
rect 876 4216 884 4224
rect 972 4216 980 4224
rect 860 4196 868 4204
rect 956 4196 964 4204
rect 892 4156 900 4164
rect 924 4156 932 4164
rect 828 4096 836 4104
rect 860 4096 868 4104
rect 668 3976 676 3984
rect 540 3816 548 3824
rect 604 3796 612 3804
rect 652 3896 660 3904
rect 636 3876 644 3884
rect 636 3856 644 3864
rect 668 3856 676 3864
rect 668 3836 676 3844
rect 636 3816 644 3824
rect 540 3776 548 3784
rect 508 3736 516 3744
rect 572 3736 580 3744
rect 700 4076 708 4084
rect 796 4036 804 4044
rect 716 4016 724 4024
rect 700 3996 708 4004
rect 700 3936 708 3944
rect 732 3936 740 3944
rect 796 3936 804 3944
rect 828 4076 836 4084
rect 844 4056 852 4064
rect 828 3916 836 3924
rect 796 3896 804 3904
rect 812 3896 820 3904
rect 700 3836 708 3844
rect 748 3836 756 3844
rect 700 3816 708 3824
rect 684 3776 692 3784
rect 652 3756 660 3764
rect 524 3656 532 3664
rect 604 3676 612 3684
rect 556 3636 564 3644
rect 572 3636 580 3644
rect 556 3576 564 3584
rect 476 3556 484 3564
rect 556 3556 564 3564
rect 572 3556 580 3564
rect 460 3536 468 3544
rect 428 3496 436 3504
rect 460 3496 468 3504
rect 428 3456 436 3464
rect 380 3416 388 3424
rect 300 3376 308 3384
rect 332 3376 340 3384
rect 412 3416 420 3424
rect 492 3476 500 3484
rect 524 3476 532 3484
rect 476 3456 484 3464
rect 460 3416 468 3424
rect 284 3356 292 3364
rect 284 3336 292 3344
rect 348 3336 356 3344
rect 252 3316 260 3324
rect 268 3276 276 3284
rect 268 3236 276 3244
rect 172 3176 180 3184
rect 172 3116 180 3124
rect 204 3116 212 3124
rect 156 3076 164 3084
rect 156 3056 164 3064
rect 12 3036 20 3044
rect 92 3036 100 3044
rect 44 3016 52 3024
rect 172 3036 180 3044
rect 188 3036 196 3044
rect 12 2896 20 2904
rect 172 2896 180 2904
rect 172 2876 180 2884
rect 92 2816 100 2824
rect 252 3036 260 3044
rect 316 3296 324 3304
rect 300 3256 308 3264
rect 316 3256 324 3264
rect 284 3196 292 3204
rect 332 3216 340 3224
rect 204 2976 212 2984
rect 220 2936 228 2944
rect 300 2956 308 2964
rect 204 2876 212 2884
rect 236 2896 244 2904
rect 236 2876 244 2884
rect 220 2816 228 2824
rect 268 2856 276 2864
rect 172 2756 180 2764
rect 108 2736 116 2744
rect 12 2696 20 2704
rect 60 2696 68 2704
rect 44 2676 52 2684
rect 92 2656 100 2664
rect 156 2696 164 2704
rect 140 2676 148 2684
rect 108 2616 116 2624
rect 284 2716 292 2724
rect 204 2696 212 2704
rect 204 2676 212 2684
rect 252 2676 260 2684
rect 316 2896 324 2904
rect 444 3376 452 3384
rect 412 3336 420 3344
rect 396 3256 404 3264
rect 412 3216 420 3224
rect 396 3196 404 3204
rect 540 3456 548 3464
rect 524 3416 532 3424
rect 492 3336 500 3344
rect 476 3276 484 3284
rect 460 3256 468 3264
rect 364 3136 372 3144
rect 380 3136 388 3144
rect 380 3056 388 3064
rect 412 3096 420 3104
rect 412 3056 420 3064
rect 380 3016 388 3024
rect 348 2956 356 2964
rect 396 2956 404 2964
rect 332 2876 340 2884
rect 316 2716 324 2724
rect 316 2696 324 2704
rect 300 2656 308 2664
rect 540 3356 548 3364
rect 492 3136 500 3144
rect 444 3116 452 3124
rect 524 3296 532 3304
rect 524 3276 532 3284
rect 524 3136 532 3144
rect 492 3096 500 3104
rect 508 3096 516 3104
rect 636 3576 644 3584
rect 652 3536 660 3544
rect 620 3516 628 3524
rect 588 3496 596 3504
rect 652 3496 660 3504
rect 764 3796 772 3804
rect 796 3796 804 3804
rect 812 3796 820 3804
rect 732 3756 740 3764
rect 780 3756 788 3764
rect 716 3716 724 3724
rect 732 3716 740 3724
rect 716 3556 724 3564
rect 604 3396 612 3404
rect 588 3356 596 3364
rect 604 3336 612 3344
rect 620 3336 628 3344
rect 604 3296 612 3304
rect 588 3276 596 3284
rect 604 3276 612 3284
rect 572 3256 580 3264
rect 556 3176 564 3184
rect 556 3096 564 3104
rect 540 3076 548 3084
rect 556 3076 564 3084
rect 492 3056 500 3064
rect 476 3036 484 3044
rect 460 2936 468 2944
rect 444 2916 452 2924
rect 428 2896 436 2904
rect 476 2896 484 2904
rect 412 2856 420 2864
rect 428 2856 436 2864
rect 364 2816 372 2824
rect 396 2776 404 2784
rect 364 2676 372 2684
rect 412 2676 420 2684
rect 252 2636 260 2644
rect 284 2636 292 2644
rect 348 2636 356 2644
rect 124 2516 132 2524
rect 12 2496 20 2504
rect 60 2496 68 2504
rect 44 2436 52 2444
rect 108 2436 116 2444
rect 12 2316 20 2324
rect 60 2396 68 2404
rect 108 2416 116 2424
rect 44 2256 52 2264
rect 92 2356 100 2364
rect 188 2536 196 2544
rect 172 2496 180 2504
rect 140 2416 148 2424
rect 140 2396 148 2404
rect 124 2356 132 2364
rect 300 2616 308 2624
rect 268 2576 276 2584
rect 236 2516 244 2524
rect 220 2496 228 2504
rect 220 2476 228 2484
rect 332 2556 340 2564
rect 316 2536 324 2544
rect 188 2396 196 2404
rect 156 2376 164 2384
rect 156 2356 164 2364
rect 204 2356 212 2364
rect 108 2276 116 2284
rect 156 2276 164 2284
rect 44 2236 52 2244
rect 12 2176 20 2184
rect 28 2136 36 2144
rect 76 2216 84 2224
rect 156 2236 164 2244
rect 92 2176 100 2184
rect 108 2176 116 2184
rect 300 2416 308 2424
rect 332 2416 340 2424
rect 316 2376 324 2384
rect 252 2356 260 2364
rect 268 2336 276 2344
rect 284 2316 292 2324
rect 412 2496 420 2504
rect 396 2456 404 2464
rect 364 2416 372 2424
rect 348 2336 356 2344
rect 380 2376 388 2384
rect 188 2296 196 2304
rect 220 2296 228 2304
rect 236 2296 244 2304
rect 348 2296 356 2304
rect 188 2216 196 2224
rect 156 2156 164 2164
rect 172 2136 180 2144
rect 108 2116 116 2124
rect 140 2116 148 2124
rect 60 2096 68 2104
rect 28 1936 36 1944
rect 76 1916 84 1924
rect 108 2056 116 2064
rect 92 1896 100 1904
rect 60 1856 68 1864
rect 12 1696 20 1704
rect 124 1936 132 1944
rect 140 1916 148 1924
rect 76 1756 84 1764
rect 60 1696 68 1704
rect 108 1696 116 1704
rect 44 1656 52 1664
rect 92 1656 100 1664
rect 92 1616 100 1624
rect 44 1596 52 1604
rect 12 1516 20 1524
rect 60 1576 68 1584
rect 12 1476 20 1484
rect 44 1316 52 1324
rect 28 1296 36 1304
rect 44 936 52 944
rect 172 1876 180 1884
rect 140 1796 148 1804
rect 252 2236 260 2244
rect 204 2196 212 2204
rect 220 2196 228 2204
rect 252 2196 260 2204
rect 204 2176 212 2184
rect 204 1956 212 1964
rect 300 2156 308 2164
rect 332 2156 340 2164
rect 236 2116 244 2124
rect 316 2116 324 2124
rect 300 2056 308 2064
rect 300 1956 308 1964
rect 220 1936 228 1944
rect 284 1936 292 1944
rect 188 1856 196 1864
rect 236 1856 244 1864
rect 268 1836 276 1844
rect 252 1816 260 1824
rect 188 1776 196 1784
rect 172 1736 180 1744
rect 236 1736 244 1744
rect 188 1716 196 1724
rect 156 1696 164 1704
rect 188 1536 196 1544
rect 124 1496 132 1504
rect 156 1496 164 1504
rect 172 1496 180 1504
rect 204 1496 212 1504
rect 156 1476 164 1484
rect 140 1416 148 1424
rect 124 1316 132 1324
rect 108 1296 116 1304
rect 220 1476 228 1484
rect 268 1616 276 1624
rect 268 1556 276 1564
rect 300 1636 308 1644
rect 332 1896 340 1904
rect 412 2336 420 2344
rect 556 3036 564 3044
rect 540 2996 548 3004
rect 588 3036 596 3044
rect 844 3836 852 3844
rect 940 4116 948 4124
rect 908 4096 916 4104
rect 908 3956 916 3964
rect 876 3936 884 3944
rect 940 3936 948 3944
rect 972 3936 980 3944
rect 892 3916 900 3924
rect 908 3916 916 3924
rect 956 3896 964 3904
rect 908 3876 916 3884
rect 940 3876 948 3884
rect 860 3816 868 3824
rect 860 3776 868 3784
rect 892 3776 900 3784
rect 828 3716 836 3724
rect 812 3696 820 3704
rect 844 3696 852 3704
rect 780 3676 788 3684
rect 908 3736 916 3744
rect 956 3816 964 3824
rect 972 3796 980 3804
rect 956 3756 964 3764
rect 940 3696 948 3704
rect 956 3696 964 3704
rect 796 3656 804 3664
rect 860 3656 868 3664
rect 956 3676 964 3684
rect 892 3636 900 3644
rect 892 3576 900 3584
rect 908 3576 916 3584
rect 924 3576 932 3584
rect 972 3576 980 3584
rect 780 3556 788 3564
rect 828 3536 836 3544
rect 860 3496 868 3504
rect 732 3456 740 3464
rect 748 3436 756 3444
rect 716 3416 724 3424
rect 748 3416 756 3424
rect 668 3396 676 3404
rect 700 3396 708 3404
rect 652 3336 660 3344
rect 700 3376 708 3384
rect 684 3356 692 3364
rect 668 3296 676 3304
rect 636 3276 644 3284
rect 620 3056 628 3064
rect 716 3276 724 3284
rect 668 3236 676 3244
rect 652 3196 660 3204
rect 652 3156 660 3164
rect 812 3476 820 3484
rect 796 3436 804 3444
rect 812 3436 820 3444
rect 876 3476 884 3484
rect 940 3536 948 3544
rect 956 3536 964 3544
rect 924 3496 932 3504
rect 844 3456 852 3464
rect 764 3276 772 3284
rect 828 3316 836 3324
rect 780 3256 788 3264
rect 732 3196 740 3204
rect 700 3136 708 3144
rect 828 3276 836 3284
rect 1004 4336 1012 4344
rect 1020 4276 1028 4284
rect 1420 4536 1428 4544
rect 1628 4536 1636 4544
rect 1116 4336 1124 4344
rect 1180 4396 1188 4404
rect 1228 4516 1236 4524
rect 1132 4316 1140 4324
rect 1132 4296 1140 4304
rect 1100 4256 1108 4264
rect 1052 4236 1060 4244
rect 1116 4236 1124 4244
rect 1036 4216 1044 4224
rect 1052 4196 1060 4204
rect 1308 4476 1316 4484
rect 1340 4496 1348 4504
rect 1420 4496 1428 4504
rect 1468 4496 1476 4504
rect 1324 4436 1332 4444
rect 1212 4376 1220 4384
rect 1260 4376 1268 4384
rect 1404 4376 1412 4384
rect 1164 4316 1172 4324
rect 1500 4496 1508 4504
rect 1740 4556 1748 4564
rect 1756 4496 1764 4504
rect 1740 4476 1748 4484
rect 1660 4436 1668 4444
rect 1566 4406 1574 4414
rect 1580 4406 1588 4414
rect 1594 4406 1602 4414
rect 1468 4376 1476 4384
rect 1484 4376 1492 4384
rect 1532 4376 1540 4384
rect 1660 4376 1668 4384
rect 1420 4356 1428 4364
rect 1340 4336 1348 4344
rect 1388 4336 1396 4344
rect 1676 4336 1684 4344
rect 1724 4336 1732 4344
rect 1420 4316 1428 4324
rect 1516 4316 1524 4324
rect 1564 4316 1572 4324
rect 1660 4316 1668 4324
rect 1692 4316 1700 4324
rect 1244 4296 1252 4304
rect 1276 4296 1284 4304
rect 1068 4176 1076 4184
rect 1404 4296 1412 4304
rect 1228 4276 1236 4284
rect 1308 4276 1316 4284
rect 1356 4276 1364 4284
rect 1276 4176 1284 4184
rect 1164 4156 1172 4164
rect 1132 4136 1140 4144
rect 1164 4136 1172 4144
rect 1036 4036 1044 4044
rect 1084 4056 1092 4064
rect 1084 4036 1092 4044
rect 1052 4016 1060 4024
rect 1036 3956 1044 3964
rect 1052 3916 1060 3924
rect 1068 3896 1076 3904
rect 1020 3876 1028 3884
rect 1020 3796 1028 3804
rect 1004 3776 1012 3784
rect 1116 4056 1124 4064
rect 1100 4016 1108 4024
rect 1100 3976 1108 3984
rect 1100 3896 1108 3904
rect 1052 3756 1060 3764
rect 1164 4116 1172 4124
rect 1212 4116 1220 4124
rect 1292 4116 1300 4124
rect 1148 3936 1156 3944
rect 1420 4236 1428 4244
rect 1324 4216 1332 4224
rect 1356 4156 1364 4164
rect 1404 4156 1412 4164
rect 1452 4296 1460 4304
rect 1500 4296 1508 4304
rect 1500 4276 1508 4284
rect 1484 4216 1492 4224
rect 1436 4196 1444 4204
rect 1532 4256 1540 4264
rect 1548 4216 1556 4224
rect 1932 4936 1940 4944
rect 1964 4936 1972 4944
rect 1836 4736 1844 4744
rect 1884 4736 1892 4744
rect 1900 4736 1908 4744
rect 1852 4696 1860 4704
rect 1900 4696 1908 4704
rect 1932 4836 1940 4844
rect 1980 4816 1988 4824
rect 1980 4796 1988 4804
rect 2028 4876 2036 4884
rect 2140 5016 2148 5024
rect 2060 4996 2068 5004
rect 2316 5036 2324 5044
rect 2188 5016 2196 5024
rect 2220 5016 2228 5024
rect 2252 5016 2260 5024
rect 2140 4936 2148 4944
rect 2044 4856 2052 4864
rect 2156 4916 2164 4924
rect 2108 4896 2116 4904
rect 2284 4976 2292 4984
rect 2332 4976 2340 4984
rect 2236 4956 2244 4964
rect 2236 4936 2244 4944
rect 2252 4916 2260 4924
rect 2300 4956 2308 4964
rect 2316 4956 2324 4964
rect 2300 4936 2308 4944
rect 2348 4936 2356 4944
rect 2124 4876 2132 4884
rect 2204 4876 2212 4884
rect 2300 4876 2308 4884
rect 2140 4816 2148 4824
rect 2124 4796 2132 4804
rect 2076 4776 2084 4784
rect 1996 4736 2004 4744
rect 1964 4696 1972 4704
rect 2028 4696 2036 4704
rect 1916 4676 1924 4684
rect 1980 4676 1988 4684
rect 1868 4656 1876 4664
rect 1932 4656 1940 4664
rect 1804 4616 1812 4624
rect 1852 4556 1860 4564
rect 1948 4556 1956 4564
rect 1932 4536 1940 4544
rect 1916 4516 1924 4524
rect 1836 4496 1844 4504
rect 1900 4496 1908 4504
rect 1804 4476 1812 4484
rect 1820 4436 1828 4444
rect 1996 4536 2004 4544
rect 1980 4516 1988 4524
rect 2028 4516 2036 4524
rect 1964 4436 1972 4444
rect 1980 4436 1988 4444
rect 1980 4376 1988 4384
rect 2012 4376 2020 4384
rect 1964 4356 1972 4364
rect 1804 4316 1812 4324
rect 1740 4296 1748 4304
rect 1708 4276 1716 4284
rect 1756 4276 1764 4284
rect 1644 4256 1652 4264
rect 1580 4196 1588 4204
rect 1868 4256 1876 4264
rect 1852 4216 1860 4224
rect 1916 4216 1924 4224
rect 1740 4196 1748 4204
rect 1996 4356 2004 4364
rect 2092 4716 2100 4724
rect 2156 4716 2164 4724
rect 2252 4716 2260 4724
rect 2220 4696 2228 4704
rect 2140 4676 2148 4684
rect 2172 4676 2180 4684
rect 2204 4656 2212 4664
rect 2140 4636 2148 4644
rect 2188 4576 2196 4584
rect 2172 4556 2180 4564
rect 2060 4536 2068 4544
rect 2108 4536 2116 4544
rect 2076 4516 2084 4524
rect 2124 4516 2132 4524
rect 2076 4496 2084 4504
rect 2060 4476 2068 4484
rect 2092 4476 2100 4484
rect 2156 4476 2164 4484
rect 2204 4456 2212 4464
rect 2092 4376 2100 4384
rect 2076 4356 2084 4364
rect 2044 4336 2052 4344
rect 2140 4336 2148 4344
rect 1964 4276 1972 4284
rect 1996 4256 2004 4264
rect 2028 4236 2036 4244
rect 2028 4216 2036 4224
rect 1708 4176 1716 4184
rect 1948 4176 1956 4184
rect 1564 4156 1572 4164
rect 1692 4156 1700 4164
rect 1356 4136 1364 4144
rect 1324 4116 1332 4124
rect 1244 4096 1252 4104
rect 1308 4096 1316 4104
rect 1356 4096 1364 4104
rect 1228 4076 1236 4084
rect 1196 4056 1204 4064
rect 1196 3956 1204 3964
rect 1180 3916 1188 3924
rect 1260 4076 1268 4084
rect 1276 3956 1284 3964
rect 1132 3876 1140 3884
rect 1164 3876 1172 3884
rect 1196 3876 1204 3884
rect 1292 3876 1300 3884
rect 1324 3876 1332 3884
rect 1340 3876 1348 3884
rect 1116 3836 1124 3844
rect 1196 3836 1204 3844
rect 1212 3836 1220 3844
rect 1212 3796 1220 3804
rect 1116 3776 1124 3784
rect 1148 3776 1156 3784
rect 1020 3696 1028 3704
rect 1068 3516 1076 3524
rect 988 3456 996 3464
rect 860 3416 868 3424
rect 940 3416 948 3424
rect 972 3416 980 3424
rect 892 3396 900 3404
rect 860 3356 868 3364
rect 876 3336 884 3344
rect 844 3216 852 3224
rect 812 3196 820 3204
rect 908 3356 916 3364
rect 860 3156 868 3164
rect 828 3136 836 3144
rect 716 3116 724 3124
rect 780 3116 788 3124
rect 700 3096 708 3104
rect 828 3096 836 3104
rect 684 3076 692 3084
rect 716 3076 724 3084
rect 812 3076 820 3084
rect 892 3096 900 3104
rect 924 3116 932 3124
rect 604 3016 612 3024
rect 572 2996 580 3004
rect 524 2956 532 2964
rect 492 2816 500 2824
rect 444 2776 452 2784
rect 476 2756 484 2764
rect 508 2736 516 2744
rect 508 2680 516 2684
rect 508 2676 516 2680
rect 460 2656 468 2664
rect 492 2656 500 2664
rect 508 2616 516 2624
rect 476 2556 484 2564
rect 508 2556 516 2564
rect 460 2536 468 2544
rect 492 2536 500 2544
rect 508 2536 516 2544
rect 556 2936 564 2944
rect 540 2896 548 2904
rect 540 2716 548 2724
rect 652 3036 660 3044
rect 588 2976 596 2984
rect 604 2916 612 2924
rect 588 2876 596 2884
rect 716 3036 724 3044
rect 748 2996 756 3004
rect 684 2976 692 2984
rect 732 2936 740 2944
rect 668 2916 676 2924
rect 636 2856 644 2864
rect 668 2856 676 2864
rect 716 2876 724 2884
rect 652 2836 660 2844
rect 684 2836 692 2844
rect 700 2836 708 2844
rect 636 2816 644 2824
rect 876 3076 884 3084
rect 860 3036 868 3044
rect 876 3036 884 3044
rect 860 3016 868 3024
rect 780 2936 788 2944
rect 860 2936 868 2944
rect 780 2916 788 2924
rect 716 2796 724 2804
rect 764 2796 772 2804
rect 700 2776 708 2784
rect 604 2716 612 2724
rect 588 2676 596 2684
rect 556 2656 564 2664
rect 620 2656 628 2664
rect 604 2616 612 2624
rect 604 2596 612 2604
rect 572 2556 580 2564
rect 444 2496 452 2504
rect 444 2336 452 2344
rect 444 2316 452 2324
rect 364 2216 372 2224
rect 380 2216 388 2224
rect 380 2116 388 2124
rect 364 1996 372 2004
rect 476 2336 484 2344
rect 460 2296 468 2304
rect 428 2116 436 2124
rect 428 1996 436 2004
rect 396 1976 404 1984
rect 508 2496 516 2504
rect 524 2436 532 2444
rect 572 2536 580 2544
rect 668 2756 676 2764
rect 652 2736 660 2744
rect 684 2716 692 2724
rect 684 2676 692 2684
rect 652 2596 660 2604
rect 652 2576 660 2584
rect 556 2496 564 2504
rect 620 2416 628 2424
rect 812 2856 820 2864
rect 908 2936 916 2944
rect 828 2836 836 2844
rect 796 2756 804 2764
rect 716 2736 724 2744
rect 764 2736 772 2744
rect 844 2736 852 2744
rect 716 2656 724 2664
rect 764 2716 772 2724
rect 796 2716 804 2724
rect 764 2656 772 2664
rect 780 2656 788 2664
rect 748 2616 756 2624
rect 812 2616 820 2624
rect 828 2616 836 2624
rect 764 2596 772 2604
rect 812 2596 820 2604
rect 828 2596 836 2604
rect 700 2556 708 2564
rect 668 2516 676 2524
rect 668 2356 676 2364
rect 636 2336 644 2344
rect 652 2336 660 2344
rect 476 2216 484 2224
rect 508 2196 516 2204
rect 508 2176 516 2184
rect 492 2156 500 2164
rect 476 2136 484 2144
rect 460 2096 468 2104
rect 508 2096 516 2104
rect 460 2056 468 2064
rect 476 2056 484 2064
rect 460 1996 468 2004
rect 380 1936 388 1944
rect 396 1896 404 1904
rect 348 1856 356 1864
rect 396 1856 404 1864
rect 348 1836 356 1844
rect 364 1836 372 1844
rect 380 1756 388 1764
rect 348 1736 356 1744
rect 364 1716 372 1724
rect 412 1716 420 1724
rect 348 1636 356 1644
rect 332 1556 340 1564
rect 412 1696 420 1704
rect 396 1596 404 1604
rect 460 1956 468 1964
rect 476 1936 484 1944
rect 668 2316 676 2324
rect 572 2296 580 2304
rect 668 2296 676 2304
rect 540 2280 548 2284
rect 540 2276 548 2280
rect 556 2256 564 2264
rect 540 2216 548 2224
rect 652 2256 660 2264
rect 588 2156 596 2164
rect 636 2156 644 2164
rect 620 2116 628 2124
rect 652 2136 660 2144
rect 604 2096 612 2104
rect 556 1996 564 2004
rect 620 1996 628 2004
rect 540 1976 548 1984
rect 524 1896 532 1904
rect 476 1876 484 1884
rect 444 1776 452 1784
rect 460 1756 468 1764
rect 444 1716 452 1724
rect 476 1676 484 1684
rect 396 1556 404 1564
rect 428 1556 436 1564
rect 412 1536 420 1544
rect 524 1816 532 1824
rect 572 1916 580 1924
rect 588 1916 596 1924
rect 588 1896 596 1904
rect 572 1756 580 1764
rect 556 1736 564 1744
rect 508 1716 516 1724
rect 556 1716 564 1724
rect 780 2536 788 2544
rect 812 2536 820 2544
rect 748 2516 756 2524
rect 876 2776 884 2784
rect 860 2696 868 2704
rect 940 3076 948 3084
rect 988 3296 996 3304
rect 1052 3476 1060 3484
rect 1100 3736 1108 3744
rect 1164 3736 1172 3744
rect 1164 3696 1172 3704
rect 1180 3636 1188 3644
rect 1132 3616 1140 3624
rect 1404 3996 1412 4004
rect 1372 3856 1380 3864
rect 1388 3856 1396 3864
rect 1420 3976 1428 3984
rect 1436 3956 1444 3964
rect 1420 3916 1428 3924
rect 1516 4076 1524 4084
rect 1884 4156 1892 4164
rect 1948 4156 1956 4164
rect 1628 4136 1636 4144
rect 1820 4136 1828 4144
rect 1468 4056 1476 4064
rect 1580 4056 1588 4064
rect 1566 4006 1574 4014
rect 1580 4006 1588 4014
rect 1594 4006 1602 4014
rect 1484 3976 1492 3984
rect 1500 3976 1508 3984
rect 1468 3936 1476 3944
rect 1452 3896 1460 3904
rect 1452 3856 1460 3864
rect 1404 3816 1412 3824
rect 1404 3796 1412 3804
rect 1372 3756 1380 3764
rect 1244 3676 1252 3684
rect 1196 3596 1204 3604
rect 1116 3496 1124 3504
rect 1100 3456 1108 3464
rect 1052 3416 1060 3424
rect 1036 3376 1044 3384
rect 1052 3356 1060 3364
rect 1036 3316 1044 3324
rect 1020 3276 1028 3284
rect 1004 3256 1012 3264
rect 1020 3216 1028 3224
rect 972 3076 980 3084
rect 1004 3076 1012 3084
rect 972 3056 980 3064
rect 1004 3056 1012 3064
rect 940 2976 948 2984
rect 956 2976 964 2984
rect 924 2896 932 2904
rect 908 2856 916 2864
rect 956 2956 964 2964
rect 956 2856 964 2864
rect 940 2836 948 2844
rect 924 2816 932 2824
rect 908 2736 916 2744
rect 1052 3196 1060 3204
rect 1052 3176 1060 3184
rect 1036 3156 1044 3164
rect 1036 3116 1044 3124
rect 1052 3096 1060 3104
rect 1036 3056 1044 3064
rect 988 2936 996 2944
rect 1084 3296 1092 3304
rect 1180 3496 1188 3504
rect 1164 3476 1172 3484
rect 1180 3476 1188 3484
rect 1148 3416 1156 3424
rect 1132 3396 1140 3404
rect 1116 3356 1124 3364
rect 1164 3356 1172 3364
rect 1132 3156 1140 3164
rect 1148 3156 1156 3164
rect 1084 3116 1092 3124
rect 1388 3716 1396 3724
rect 1308 3636 1316 3644
rect 1276 3596 1284 3604
rect 1276 3576 1284 3584
rect 1260 3556 1268 3564
rect 1244 3536 1252 3544
rect 1212 3516 1220 3524
rect 1228 3516 1236 3524
rect 1212 3436 1220 3444
rect 1292 3556 1300 3564
rect 1340 3556 1348 3564
rect 1308 3536 1316 3544
rect 1356 3536 1364 3544
rect 1516 3876 1524 3884
rect 1612 3876 1620 3884
rect 1676 4116 1684 4124
rect 1660 4076 1668 4084
rect 1644 3976 1652 3984
rect 2012 4136 2020 4144
rect 1868 4116 1876 4124
rect 1916 4116 1924 4124
rect 1996 4116 2004 4124
rect 1836 4076 1844 4084
rect 1980 4076 1988 4084
rect 1804 4056 1812 4064
rect 1836 4016 1844 4024
rect 1964 3996 1972 4004
rect 1996 3996 2004 4004
rect 2092 4216 2100 4224
rect 2108 4196 2116 4204
rect 2044 4176 2052 4184
rect 2108 4156 2116 4164
rect 2044 4136 2052 4144
rect 2060 4116 2068 4124
rect 2076 4116 2084 4124
rect 2108 4056 2116 4064
rect 2076 4036 2084 4044
rect 2124 4036 2132 4044
rect 2028 3996 2036 4004
rect 1916 3956 1924 3964
rect 1900 3916 1908 3924
rect 2044 3916 2052 3924
rect 1660 3896 1668 3904
rect 1868 3896 1876 3904
rect 1964 3896 1972 3904
rect 1996 3896 2004 3904
rect 1580 3816 1588 3824
rect 1484 3796 1492 3804
rect 1436 3756 1444 3764
rect 1548 3736 1556 3744
rect 1436 3716 1444 3724
rect 1452 3716 1460 3724
rect 1532 3716 1540 3724
rect 1548 3716 1556 3724
rect 1740 3836 1748 3844
rect 1628 3816 1636 3824
rect 1708 3816 1716 3824
rect 1708 3776 1716 3784
rect 1788 3816 1796 3824
rect 1772 3796 1780 3804
rect 1500 3696 1508 3704
rect 1612 3696 1620 3704
rect 1420 3676 1428 3684
rect 1436 3676 1444 3684
rect 1468 3656 1476 3664
rect 1436 3636 1444 3644
rect 1452 3636 1460 3644
rect 1404 3516 1412 3524
rect 1420 3516 1428 3524
rect 1566 3606 1574 3614
rect 1580 3606 1588 3614
rect 1594 3606 1602 3614
rect 1532 3596 1540 3604
rect 1500 3556 1508 3564
rect 1532 3556 1540 3564
rect 1308 3496 1316 3504
rect 1356 3496 1364 3504
rect 1388 3496 1396 3504
rect 1436 3496 1444 3504
rect 1420 3456 1428 3464
rect 1276 3416 1284 3424
rect 1308 3416 1316 3424
rect 1340 3416 1348 3424
rect 1372 3416 1380 3424
rect 1276 3396 1284 3404
rect 1388 3396 1396 3404
rect 1308 3376 1316 3384
rect 1324 3376 1332 3384
rect 1372 3356 1380 3364
rect 1180 3276 1188 3284
rect 1180 3196 1188 3204
rect 1084 3076 1092 3084
rect 1116 3096 1124 3104
rect 1068 2876 1076 2884
rect 1020 2856 1028 2864
rect 1036 2796 1044 2804
rect 1116 2936 1124 2944
rect 1100 2856 1108 2864
rect 1164 3116 1172 3124
rect 1180 3096 1188 3104
rect 1484 3476 1492 3484
rect 1564 3536 1572 3544
rect 1612 3536 1620 3544
rect 1820 3856 1828 3864
rect 1836 3856 1844 3864
rect 1868 3856 1876 3864
rect 1884 3856 1892 3864
rect 1932 3856 1940 3864
rect 1980 3856 1988 3864
rect 1820 3816 1828 3824
rect 1756 3716 1764 3724
rect 1772 3716 1780 3724
rect 1676 3696 1684 3704
rect 1644 3676 1652 3684
rect 1660 3656 1668 3664
rect 1644 3556 1652 3564
rect 1580 3516 1588 3524
rect 1628 3516 1636 3524
rect 1596 3496 1604 3504
rect 1580 3476 1588 3484
rect 1596 3436 1604 3444
rect 1580 3416 1588 3424
rect 1468 3396 1476 3404
rect 1516 3396 1524 3404
rect 1244 3336 1252 3344
rect 1292 3336 1300 3344
rect 1340 3316 1348 3324
rect 1404 3316 1412 3324
rect 1276 3296 1284 3304
rect 1324 3296 1332 3304
rect 1372 3276 1380 3284
rect 1244 3236 1252 3244
rect 1292 3236 1300 3244
rect 1228 3216 1236 3224
rect 1228 3116 1236 3124
rect 1244 3096 1252 3104
rect 1212 3016 1220 3024
rect 1196 2996 1204 3004
rect 1164 2976 1172 2984
rect 1276 3176 1284 3184
rect 1276 3056 1284 3064
rect 1340 3156 1348 3164
rect 1308 3136 1316 3144
rect 1324 3136 1332 3144
rect 1452 3356 1460 3364
rect 1436 3336 1444 3344
rect 1548 3336 1556 3344
rect 1436 3296 1444 3304
rect 1612 3416 1620 3424
rect 1660 3416 1668 3424
rect 1852 3836 1860 3844
rect 1852 3776 1860 3784
rect 1884 3776 1892 3784
rect 2060 3876 2068 3884
rect 2188 4316 2196 4324
rect 2204 4256 2212 4264
rect 2284 4576 2292 4584
rect 2268 4556 2276 4564
rect 2268 4516 2276 4524
rect 2252 4436 2260 4444
rect 2268 4416 2276 4424
rect 2428 5076 2436 5084
rect 2412 5036 2420 5044
rect 2428 5036 2436 5044
rect 2572 5076 2580 5084
rect 2572 5056 2580 5064
rect 2524 5016 2532 5024
rect 2412 4996 2420 5004
rect 2476 4996 2484 5004
rect 2380 4956 2388 4964
rect 2380 4936 2388 4944
rect 2460 4956 2468 4964
rect 2444 4896 2452 4904
rect 2428 4876 2436 4884
rect 2364 4836 2372 4844
rect 2428 4756 2436 4764
rect 2508 4976 2516 4984
rect 2524 4956 2532 4964
rect 2524 4896 2532 4904
rect 2588 5036 2596 5044
rect 2668 5076 2676 5084
rect 2620 5056 2628 5064
rect 2652 5056 2660 5064
rect 2732 5076 2740 5084
rect 2828 5096 2836 5104
rect 2892 5096 2900 5104
rect 2988 5096 2996 5104
rect 2956 5076 2964 5084
rect 2700 5056 2708 5064
rect 2764 5056 2772 5064
rect 2908 5056 2916 5064
rect 2684 5036 2692 5044
rect 2604 4996 2612 5004
rect 2556 4976 2564 4984
rect 2620 4956 2628 4964
rect 2668 4956 2676 4964
rect 2732 4956 2740 4964
rect 2572 4936 2580 4944
rect 2860 4976 2868 4984
rect 2924 4976 2932 4984
rect 2636 4936 2644 4944
rect 2796 4936 2804 4944
rect 2556 4916 2564 4924
rect 2588 4916 2596 4924
rect 2652 4916 2660 4924
rect 2572 4896 2580 4904
rect 2620 4896 2628 4904
rect 2492 4876 2500 4884
rect 2700 4876 2708 4884
rect 2716 4876 2724 4884
rect 2460 4736 2468 4744
rect 2476 4716 2484 4724
rect 2460 4696 2468 4704
rect 2348 4656 2356 4664
rect 2332 4556 2340 4564
rect 2316 4536 2324 4544
rect 2428 4656 2436 4664
rect 2364 4636 2372 4644
rect 2396 4556 2404 4564
rect 2412 4556 2420 4564
rect 2444 4636 2452 4644
rect 2412 4536 2420 4544
rect 2460 4616 2468 4624
rect 2524 4776 2532 4784
rect 2572 4756 2580 4764
rect 2508 4736 2516 4744
rect 2700 4776 2708 4784
rect 2652 4756 2660 4764
rect 2588 4736 2596 4744
rect 2620 4736 2628 4744
rect 2556 4716 2564 4724
rect 2572 4716 2580 4724
rect 2652 4716 2660 4724
rect 2492 4696 2500 4704
rect 2524 4696 2532 4704
rect 2604 4696 2612 4704
rect 2844 4896 2852 4904
rect 2956 4996 2964 5004
rect 2940 4936 2948 4944
rect 2908 4916 2916 4924
rect 2940 4896 2948 4904
rect 2876 4876 2884 4884
rect 2812 4856 2820 4864
rect 2732 4716 2740 4724
rect 2764 4716 2772 4724
rect 2716 4696 2724 4704
rect 2540 4676 2548 4684
rect 2668 4676 2676 4684
rect 2636 4656 2644 4664
rect 2348 4396 2356 4404
rect 2284 4316 2292 4324
rect 2300 4316 2308 4324
rect 2268 4296 2276 4304
rect 2220 4196 2228 4204
rect 2156 4136 2164 4144
rect 2156 4116 2164 4124
rect 2236 4136 2244 4144
rect 2268 4236 2276 4244
rect 2268 4176 2276 4184
rect 2252 4116 2260 4124
rect 2204 4076 2212 4084
rect 2188 4056 2196 4064
rect 2156 4036 2164 4044
rect 2140 3936 2148 3944
rect 2252 4076 2260 4084
rect 2236 4056 2244 4064
rect 2668 4616 2676 4624
rect 2700 4616 2708 4624
rect 2620 4576 2628 4584
rect 2492 4556 2500 4564
rect 2588 4556 2596 4564
rect 2668 4556 2676 4564
rect 2540 4516 2548 4524
rect 2572 4516 2580 4524
rect 2476 4496 2484 4504
rect 2524 4496 2532 4504
rect 2556 4496 2564 4504
rect 2652 4516 2660 4524
rect 2652 4476 2660 4484
rect 2492 4456 2500 4464
rect 2508 4456 2516 4464
rect 2492 4436 2500 4444
rect 2460 4396 2468 4404
rect 2396 4376 2404 4384
rect 2428 4336 2436 4344
rect 2396 4316 2404 4324
rect 2444 4316 2452 4324
rect 2300 4256 2308 4264
rect 2284 4136 2292 4144
rect 2396 4296 2404 4304
rect 2364 4276 2372 4284
rect 2412 4276 2420 4284
rect 2332 4236 2340 4244
rect 2364 4216 2372 4224
rect 2380 4176 2388 4184
rect 2412 4156 2420 4164
rect 2460 4276 2468 4284
rect 2460 4196 2468 4204
rect 2316 4136 2324 4144
rect 2396 4136 2404 4144
rect 2300 4116 2308 4124
rect 2428 4116 2436 4124
rect 2476 4156 2484 4164
rect 2316 4096 2324 4104
rect 2268 4036 2276 4044
rect 2220 4016 2228 4024
rect 2220 3996 2228 4004
rect 2236 3976 2244 3984
rect 2204 3956 2212 3964
rect 2252 3876 2260 3884
rect 2172 3836 2180 3844
rect 2124 3796 2132 3804
rect 1932 3756 1940 3764
rect 1996 3756 2004 3764
rect 2044 3756 2052 3764
rect 1980 3736 1988 3744
rect 2060 3736 2068 3744
rect 2092 3736 2100 3744
rect 1820 3716 1828 3724
rect 1868 3716 1876 3724
rect 1948 3716 1956 3724
rect 2012 3716 2020 3724
rect 2092 3716 2100 3724
rect 2188 3796 2196 3804
rect 2140 3716 2148 3724
rect 2204 3716 2212 3724
rect 1804 3636 1812 3644
rect 1884 3636 1892 3644
rect 1932 3636 1940 3644
rect 1708 3596 1716 3604
rect 1788 3596 1796 3604
rect 1692 3516 1700 3524
rect 1740 3556 1748 3564
rect 1804 3556 1812 3564
rect 1788 3516 1796 3524
rect 2108 3676 2116 3684
rect 2044 3656 2052 3664
rect 2012 3596 2020 3604
rect 1980 3576 1988 3584
rect 1964 3516 1972 3524
rect 1852 3496 1860 3504
rect 1740 3476 1748 3484
rect 1772 3476 1780 3484
rect 1948 3476 1956 3484
rect 1980 3476 1988 3484
rect 1692 3456 1700 3464
rect 1708 3456 1716 3464
rect 1772 3456 1780 3464
rect 1788 3456 1796 3464
rect 1596 3376 1604 3384
rect 1676 3376 1684 3384
rect 1612 3356 1620 3364
rect 1676 3356 1684 3364
rect 1644 3336 1652 3344
rect 1644 3316 1652 3324
rect 1852 3436 1860 3444
rect 1868 3436 1876 3444
rect 1724 3336 1732 3344
rect 1788 3336 1796 3344
rect 1740 3316 1748 3324
rect 1804 3316 1812 3324
rect 1580 3256 1588 3264
rect 1804 3276 1812 3284
rect 1772 3236 1780 3244
rect 1566 3206 1574 3214
rect 1580 3206 1588 3214
rect 1594 3206 1602 3214
rect 1500 3176 1508 3184
rect 1532 3176 1540 3184
rect 1452 3156 1460 3164
rect 1372 3136 1380 3144
rect 1388 3136 1396 3144
rect 1420 3136 1428 3144
rect 1324 3116 1332 3124
rect 1308 3096 1316 3104
rect 1228 2916 1236 2924
rect 1260 2916 1268 2924
rect 1148 2896 1156 2904
rect 1228 2896 1236 2904
rect 1100 2796 1108 2804
rect 1036 2756 1044 2764
rect 1084 2756 1092 2764
rect 1004 2736 1012 2744
rect 972 2696 980 2704
rect 1004 2696 1012 2704
rect 908 2656 916 2664
rect 924 2656 932 2664
rect 988 2656 996 2664
rect 892 2636 900 2644
rect 924 2636 932 2644
rect 876 2596 884 2604
rect 892 2596 900 2604
rect 812 2476 820 2484
rect 748 2456 756 2464
rect 860 2476 868 2484
rect 844 2436 852 2444
rect 748 2316 756 2324
rect 828 2316 836 2324
rect 860 2316 868 2324
rect 956 2616 964 2624
rect 1020 2616 1028 2624
rect 1052 2716 1060 2724
rect 1052 2676 1060 2684
rect 1068 2656 1076 2664
rect 1068 2596 1076 2604
rect 1052 2556 1060 2564
rect 908 2456 916 2464
rect 924 2456 932 2464
rect 1004 2456 1012 2464
rect 1036 2436 1044 2444
rect 956 2396 964 2404
rect 700 2296 708 2304
rect 716 2296 724 2304
rect 828 2296 836 2304
rect 892 2296 900 2304
rect 908 2296 916 2304
rect 940 2296 948 2304
rect 700 2276 708 2284
rect 764 2256 772 2264
rect 796 2236 804 2244
rect 748 2196 756 2204
rect 684 2156 692 2164
rect 700 2116 708 2124
rect 700 2096 708 2104
rect 684 2076 692 2084
rect 636 1896 644 1904
rect 604 1756 612 1764
rect 524 1696 532 1704
rect 588 1696 596 1704
rect 492 1636 500 1644
rect 508 1636 516 1644
rect 428 1516 436 1524
rect 476 1516 484 1524
rect 364 1496 372 1504
rect 396 1496 404 1504
rect 284 1476 292 1484
rect 316 1476 324 1484
rect 204 1456 212 1464
rect 284 1456 292 1464
rect 220 1376 228 1384
rect 204 1336 212 1344
rect 140 1276 148 1284
rect 172 1276 180 1284
rect 172 1256 180 1264
rect 108 1116 116 1124
rect 92 1096 100 1104
rect 108 1076 116 1084
rect 156 1096 164 1104
rect 156 1056 164 1064
rect 124 976 132 984
rect 92 956 100 964
rect 108 936 116 944
rect 76 916 84 924
rect 140 956 148 964
rect 28 876 36 884
rect 124 896 132 904
rect 140 896 148 904
rect 76 876 84 884
rect 60 716 68 724
rect 76 696 84 704
rect 92 676 100 684
rect 60 636 68 644
rect 252 1376 260 1384
rect 236 1356 244 1364
rect 236 1336 244 1344
rect 316 1376 324 1384
rect 268 1296 276 1304
rect 188 1116 196 1124
rect 204 1116 212 1124
rect 284 1276 292 1284
rect 460 1476 468 1484
rect 508 1476 516 1484
rect 348 1416 356 1424
rect 348 1376 356 1384
rect 332 1296 340 1304
rect 348 1276 356 1284
rect 300 1236 308 1244
rect 268 1116 276 1124
rect 220 1096 228 1104
rect 204 1076 212 1084
rect 188 1056 196 1064
rect 204 956 212 964
rect 188 936 196 944
rect 220 936 228 944
rect 236 936 244 944
rect 284 956 292 964
rect 412 1356 420 1364
rect 396 1296 404 1304
rect 556 1536 564 1544
rect 524 1416 532 1424
rect 492 1396 500 1404
rect 524 1396 532 1404
rect 492 1356 500 1364
rect 476 1336 484 1344
rect 460 1296 468 1304
rect 380 1276 388 1284
rect 444 1276 452 1284
rect 364 1256 372 1264
rect 492 1236 500 1244
rect 348 1196 356 1204
rect 316 1116 324 1124
rect 348 1116 356 1124
rect 396 1196 404 1204
rect 588 1616 596 1624
rect 588 1516 596 1524
rect 572 1476 580 1484
rect 636 1796 644 1804
rect 636 1716 644 1724
rect 620 1576 628 1584
rect 668 1916 676 1924
rect 780 2116 788 2124
rect 924 2256 932 2264
rect 988 2316 996 2324
rect 1020 2296 1028 2304
rect 1036 2296 1044 2304
rect 1036 2256 1044 2264
rect 828 2236 836 2244
rect 844 2196 852 2204
rect 860 2196 868 2204
rect 876 2176 884 2184
rect 908 2156 916 2164
rect 876 2136 884 2144
rect 956 2236 964 2244
rect 956 2216 964 2224
rect 1036 2196 1044 2204
rect 1004 2156 1012 2164
rect 972 2136 980 2144
rect 716 2056 724 2064
rect 780 2056 788 2064
rect 732 2036 740 2044
rect 748 2036 756 2044
rect 748 1956 756 1964
rect 876 1996 884 2004
rect 1020 2136 1028 2144
rect 1036 2136 1044 2144
rect 1100 2616 1108 2624
rect 1100 2556 1108 2564
rect 1084 2496 1092 2504
rect 1100 2496 1108 2504
rect 1068 2436 1076 2444
rect 1068 2316 1076 2324
rect 1100 2316 1108 2324
rect 1084 2296 1092 2304
rect 1132 2796 1140 2804
rect 1260 2796 1268 2804
rect 1244 2776 1252 2784
rect 1180 2736 1188 2744
rect 1164 2716 1172 2724
rect 1212 2696 1220 2704
rect 1228 2696 1236 2704
rect 1148 2656 1156 2664
rect 1228 2656 1236 2664
rect 1164 2596 1172 2604
rect 1148 2556 1156 2564
rect 1132 2536 1140 2544
rect 1340 3076 1348 3084
rect 1324 3016 1332 3024
rect 1420 3116 1428 3124
rect 1468 3096 1476 3104
rect 1548 3156 1556 3164
rect 1628 3156 1636 3164
rect 1516 3136 1524 3144
rect 1564 3096 1572 3104
rect 1676 3116 1684 3124
rect 1660 3096 1668 3104
rect 1804 3216 1812 3224
rect 1932 3396 1940 3404
rect 1980 3356 1988 3364
rect 1916 3316 1924 3324
rect 2188 3556 2196 3564
rect 2236 3556 2244 3564
rect 2188 3536 2196 3544
rect 2076 3516 2084 3524
rect 2028 3476 2036 3484
rect 2092 3476 2100 3484
rect 2140 3476 2148 3484
rect 2172 3516 2180 3524
rect 2156 3416 2164 3424
rect 2156 3336 2164 3344
rect 2044 3316 2052 3324
rect 2092 3316 2100 3324
rect 2124 3316 2132 3324
rect 1884 3296 1892 3304
rect 1964 3296 1972 3304
rect 1868 3236 1876 3244
rect 1964 3236 1972 3244
rect 1852 3156 1860 3164
rect 1772 3136 1780 3144
rect 1836 3136 1844 3144
rect 2012 3196 2020 3204
rect 1996 3156 2004 3164
rect 1948 3136 1956 3144
rect 1996 3136 2004 3144
rect 2060 3276 2068 3284
rect 2076 3156 2084 3164
rect 2124 3296 2132 3304
rect 2108 3276 2116 3284
rect 2204 3496 2212 3504
rect 2220 3476 2228 3484
rect 2268 3856 2276 3864
rect 2300 3836 2308 3844
rect 2284 3756 2292 3764
rect 2268 3716 2276 3724
rect 2268 3676 2276 3684
rect 2460 4056 2468 4064
rect 2332 4036 2340 4044
rect 2332 3936 2340 3944
rect 2716 4456 2724 4464
rect 2684 4416 2692 4424
rect 2716 4416 2724 4424
rect 2572 4356 2580 4364
rect 2508 4336 2516 4344
rect 2588 4336 2596 4344
rect 2636 4336 2644 4344
rect 2668 4336 2676 4344
rect 2556 4296 2564 4304
rect 2796 4696 2804 4704
rect 2860 4756 2868 4764
rect 2844 4736 2852 4744
rect 2748 4456 2756 4464
rect 2748 4436 2756 4444
rect 2732 4316 2740 4324
rect 2796 4656 2804 4664
rect 2828 4656 2836 4664
rect 2828 4596 2836 4604
rect 2780 4536 2788 4544
rect 2812 4516 2820 4524
rect 2780 4496 2788 4504
rect 2812 4496 2820 4504
rect 2604 4296 2612 4304
rect 2748 4296 2756 4304
rect 2732 4276 2740 4284
rect 2764 4276 2772 4284
rect 2540 4256 2548 4264
rect 2620 4256 2628 4264
rect 2684 4256 2692 4264
rect 2572 4196 2580 4204
rect 2540 4176 2548 4184
rect 2556 4176 2564 4184
rect 2508 4136 2516 4144
rect 2348 3756 2356 3764
rect 2396 3876 2404 3884
rect 2380 3856 2388 3864
rect 2396 3816 2404 3824
rect 2380 3796 2388 3804
rect 2332 3696 2340 3704
rect 2364 3696 2372 3704
rect 2316 3676 2324 3684
rect 2396 3676 2404 3684
rect 2380 3636 2388 3644
rect 2364 3616 2372 3624
rect 2348 3596 2356 3604
rect 2300 3576 2308 3584
rect 2284 3536 2292 3544
rect 2348 3536 2356 3544
rect 2300 3496 2308 3504
rect 2332 3496 2340 3504
rect 2300 3476 2308 3484
rect 2364 3496 2372 3504
rect 2348 3476 2356 3484
rect 2268 3436 2276 3444
rect 2188 3396 2196 3404
rect 2236 3396 2244 3404
rect 2332 3416 2340 3424
rect 2364 3416 2372 3424
rect 2316 3396 2324 3404
rect 2300 3376 2308 3384
rect 2284 3336 2292 3344
rect 2220 3316 2228 3324
rect 2188 3296 2196 3304
rect 2172 3236 2180 3244
rect 2124 3156 2132 3164
rect 2108 3136 2116 3144
rect 1868 3116 1876 3124
rect 1740 3096 1748 3104
rect 1724 3076 1732 3084
rect 1356 3056 1364 3064
rect 1388 3056 1396 3064
rect 1452 3056 1460 3064
rect 1500 3056 1508 3064
rect 1516 3056 1524 3064
rect 1388 2996 1396 3004
rect 1372 2976 1380 2984
rect 1388 2916 1396 2924
rect 1420 3036 1428 3044
rect 1756 3036 1764 3044
rect 1676 3016 1684 3024
rect 1484 2976 1492 2984
rect 1452 2956 1460 2964
rect 1436 2936 1444 2944
rect 1404 2896 1412 2904
rect 1324 2856 1332 2864
rect 1388 2796 1396 2804
rect 1372 2696 1380 2704
rect 1276 2616 1284 2624
rect 1164 2496 1172 2504
rect 1132 2476 1140 2484
rect 1244 2576 1252 2584
rect 1356 2656 1364 2664
rect 1420 2776 1428 2784
rect 1404 2736 1412 2744
rect 1420 2736 1428 2744
rect 1516 2996 1524 3004
rect 1580 2996 1588 3004
rect 1612 2996 1620 3004
rect 1692 2976 1700 2984
rect 2012 3096 2020 3104
rect 1852 3076 1860 3084
rect 1804 3056 1812 3064
rect 1836 3056 1844 3064
rect 1932 3076 1940 3084
rect 2012 3076 2020 3084
rect 2076 3096 2084 3104
rect 2204 3276 2212 3284
rect 2268 3256 2276 3264
rect 2204 3176 2212 3184
rect 2252 3176 2260 3184
rect 2140 3116 2148 3124
rect 2172 3116 2180 3124
rect 2188 3116 2196 3124
rect 2220 3116 2228 3124
rect 2188 3076 2196 3084
rect 1868 3036 1876 3044
rect 1916 3036 1924 3044
rect 1884 2996 1892 3004
rect 1932 2996 1940 3004
rect 1788 2956 1796 2964
rect 1804 2956 1812 2964
rect 1852 2956 1860 2964
rect 1532 2936 1540 2944
rect 1644 2936 1652 2944
rect 1740 2936 1748 2944
rect 1788 2936 1796 2944
rect 1468 2916 1476 2924
rect 1708 2916 1716 2924
rect 1772 2916 1780 2924
rect 1452 2896 1460 2904
rect 1628 2896 1636 2904
rect 1566 2806 1574 2814
rect 1580 2806 1588 2814
rect 1594 2806 1602 2814
rect 1500 2796 1508 2804
rect 1468 2736 1476 2744
rect 1484 2676 1492 2684
rect 1388 2636 1396 2644
rect 1388 2616 1396 2624
rect 1404 2616 1412 2624
rect 1452 2616 1460 2624
rect 1340 2596 1348 2604
rect 1404 2596 1412 2604
rect 1292 2536 1300 2544
rect 1276 2516 1284 2524
rect 1228 2496 1236 2504
rect 1180 2416 1188 2424
rect 1228 2416 1236 2424
rect 1116 2276 1124 2284
rect 1148 2276 1156 2284
rect 1068 2236 1076 2244
rect 1084 2236 1092 2244
rect 1068 2196 1076 2204
rect 1212 2316 1220 2324
rect 1196 2296 1204 2304
rect 1180 2256 1188 2264
rect 1196 2236 1204 2244
rect 1116 2176 1124 2184
rect 1212 2176 1220 2184
rect 1356 2476 1364 2484
rect 1436 2576 1444 2584
rect 1420 2476 1428 2484
rect 1404 2456 1412 2464
rect 1324 2416 1332 2424
rect 1276 2316 1284 2324
rect 1308 2316 1316 2324
rect 1292 2296 1300 2304
rect 1244 2256 1252 2264
rect 1244 2196 1252 2204
rect 1068 2136 1076 2144
rect 1180 2136 1188 2144
rect 1052 2116 1060 2124
rect 988 2056 996 2064
rect 1036 2056 1044 2064
rect 1180 2096 1188 2104
rect 940 2036 948 2044
rect 812 1936 820 1944
rect 796 1916 804 1924
rect 892 1916 900 1924
rect 684 1876 692 1884
rect 684 1816 692 1824
rect 668 1776 676 1784
rect 732 1896 740 1904
rect 812 1896 820 1904
rect 876 1896 884 1904
rect 860 1876 868 1884
rect 732 1856 740 1864
rect 716 1796 724 1804
rect 716 1776 724 1784
rect 700 1756 708 1764
rect 700 1736 708 1744
rect 860 1856 868 1864
rect 764 1836 772 1844
rect 748 1796 756 1804
rect 748 1756 756 1764
rect 764 1756 772 1764
rect 716 1716 724 1724
rect 716 1636 724 1644
rect 796 1776 804 1784
rect 796 1736 804 1744
rect 780 1636 788 1644
rect 668 1596 676 1604
rect 732 1596 740 1604
rect 844 1816 852 1824
rect 828 1756 836 1764
rect 1020 1996 1028 2004
rect 1052 1996 1060 2004
rect 956 1976 964 1984
rect 972 1976 980 1984
rect 956 1916 964 1924
rect 1004 1916 1012 1924
rect 940 1896 948 1904
rect 1004 1896 1012 1904
rect 1100 2056 1108 2064
rect 1084 2036 1092 2044
rect 1036 1916 1044 1924
rect 940 1876 948 1884
rect 956 1876 964 1884
rect 1020 1876 1028 1884
rect 908 1856 916 1864
rect 1020 1856 1028 1864
rect 924 1816 932 1824
rect 940 1756 948 1764
rect 1036 1796 1044 1804
rect 1068 1916 1076 1924
rect 1068 1816 1076 1824
rect 1068 1776 1076 1784
rect 892 1736 900 1744
rect 924 1736 932 1744
rect 956 1716 964 1724
rect 860 1676 868 1684
rect 876 1656 884 1664
rect 892 1656 900 1664
rect 844 1576 852 1584
rect 652 1536 660 1544
rect 668 1516 676 1524
rect 812 1536 820 1544
rect 620 1496 628 1504
rect 652 1496 660 1504
rect 604 1456 612 1464
rect 588 1436 596 1444
rect 604 1416 612 1424
rect 556 1396 564 1404
rect 636 1376 644 1384
rect 620 1356 628 1364
rect 684 1476 692 1484
rect 876 1616 884 1624
rect 1100 2016 1108 2024
rect 1116 2016 1124 2024
rect 1148 1996 1156 2004
rect 1132 1936 1140 1944
rect 1100 1916 1108 1924
rect 1228 1996 1236 2004
rect 1180 1956 1188 1964
rect 1212 1956 1220 1964
rect 1164 1936 1172 1944
rect 1116 1896 1124 1904
rect 1148 1896 1156 1904
rect 1116 1856 1124 1864
rect 1148 1856 1156 1864
rect 1004 1716 1012 1724
rect 1036 1716 1044 1724
rect 1084 1716 1092 1724
rect 1020 1676 1028 1684
rect 1004 1656 1012 1664
rect 924 1576 932 1584
rect 972 1576 980 1584
rect 988 1576 996 1584
rect 860 1516 868 1524
rect 908 1536 916 1544
rect 700 1456 708 1464
rect 844 1476 852 1484
rect 892 1476 900 1484
rect 732 1456 740 1464
rect 764 1456 772 1464
rect 796 1456 804 1464
rect 860 1456 868 1464
rect 716 1436 724 1444
rect 668 1356 676 1364
rect 636 1336 644 1344
rect 716 1336 724 1344
rect 540 1136 548 1144
rect 332 976 340 984
rect 380 956 388 964
rect 348 936 356 944
rect 332 916 340 924
rect 524 1096 532 1104
rect 620 1156 628 1164
rect 572 1116 580 1124
rect 684 1316 692 1324
rect 700 1296 708 1304
rect 748 1436 756 1444
rect 748 1396 756 1404
rect 748 1356 756 1364
rect 748 1336 756 1344
rect 844 1436 852 1444
rect 828 1416 836 1424
rect 780 1356 788 1364
rect 812 1336 820 1344
rect 780 1296 788 1304
rect 812 1296 820 1304
rect 732 1256 740 1264
rect 684 1236 692 1244
rect 684 1196 692 1204
rect 588 1096 596 1104
rect 636 1096 644 1104
rect 652 1096 660 1104
rect 716 1176 724 1184
rect 764 1176 772 1184
rect 796 1176 804 1184
rect 700 1156 708 1164
rect 444 1076 452 1084
rect 508 1076 516 1084
rect 572 1076 580 1084
rect 652 1076 660 1084
rect 668 1076 676 1084
rect 412 1056 420 1064
rect 524 1036 532 1044
rect 668 1036 676 1044
rect 428 996 436 1004
rect 428 956 436 964
rect 492 956 500 964
rect 412 916 420 924
rect 476 916 484 924
rect 444 896 452 904
rect 540 996 548 1004
rect 620 996 628 1004
rect 700 956 708 964
rect 700 936 708 944
rect 732 1156 740 1164
rect 748 1056 756 1064
rect 892 1416 900 1424
rect 876 1396 884 1404
rect 956 1516 964 1524
rect 924 1476 932 1484
rect 924 1396 932 1404
rect 908 1376 916 1384
rect 924 1376 932 1384
rect 924 1316 932 1324
rect 1036 1556 1044 1564
rect 1212 1936 1220 1944
rect 1196 1896 1204 1904
rect 1196 1796 1204 1804
rect 1228 1796 1236 1804
rect 1196 1756 1204 1764
rect 1212 1756 1220 1764
rect 1276 2196 1284 2204
rect 1260 2116 1268 2124
rect 1420 2396 1428 2404
rect 1532 2776 1540 2784
rect 1564 2776 1572 2784
rect 1516 2716 1524 2724
rect 1548 2676 1556 2684
rect 1500 2616 1508 2624
rect 1532 2616 1540 2624
rect 1484 2576 1492 2584
rect 1516 2576 1524 2584
rect 1468 2516 1476 2524
rect 1484 2516 1492 2524
rect 1452 2416 1460 2424
rect 1468 2376 1476 2384
rect 1372 2316 1380 2324
rect 1340 2296 1348 2304
rect 1436 2316 1444 2324
rect 1452 2296 1460 2304
rect 1692 2876 1700 2884
rect 1676 2856 1684 2864
rect 1644 2756 1652 2764
rect 1676 2716 1684 2724
rect 1804 2896 1812 2904
rect 2236 3056 2244 3064
rect 1996 3036 2004 3044
rect 2044 3036 2052 3044
rect 2108 3036 2116 3044
rect 1964 2996 1972 3004
rect 1948 2976 1956 2984
rect 1868 2916 1876 2924
rect 1884 2916 1892 2924
rect 1836 2896 1844 2904
rect 1740 2876 1748 2884
rect 1788 2876 1796 2884
rect 1724 2856 1732 2864
rect 1724 2836 1732 2844
rect 1932 2876 1940 2884
rect 1980 2916 1988 2924
rect 2012 3016 2020 3024
rect 2060 2976 2068 2984
rect 2092 2976 2100 2984
rect 2044 2956 2052 2964
rect 2028 2936 2036 2944
rect 2012 2916 2020 2924
rect 1996 2896 2004 2904
rect 2204 2996 2212 3004
rect 2364 3356 2372 3364
rect 2380 3296 2388 3304
rect 2348 3276 2356 3284
rect 2332 3216 2340 3224
rect 2316 3196 2324 3204
rect 2348 3196 2356 3204
rect 2556 4156 2564 4164
rect 2572 4096 2580 4104
rect 2732 4196 2740 4204
rect 2700 4156 2708 4164
rect 2748 4176 2756 4184
rect 2652 4116 2660 4124
rect 2684 4116 2692 4124
rect 2652 4096 2660 4104
rect 2636 4076 2644 4084
rect 2636 4036 2644 4044
rect 2652 4036 2660 4044
rect 2556 3936 2564 3944
rect 2604 3936 2612 3944
rect 2540 3916 2548 3924
rect 2572 3916 2580 3924
rect 2620 3916 2628 3924
rect 2508 3856 2516 3864
rect 2588 3836 2596 3844
rect 2508 3816 2516 3824
rect 2572 3796 2580 3804
rect 2492 3776 2500 3784
rect 2476 3756 2484 3764
rect 2508 3756 2516 3764
rect 2508 3736 2516 3744
rect 2572 3736 2580 3744
rect 2444 3716 2452 3724
rect 2460 3716 2468 3724
rect 2492 3696 2500 3704
rect 2524 3676 2532 3684
rect 2412 3656 2420 3664
rect 2428 3616 2436 3624
rect 2524 3636 2532 3644
rect 2508 3576 2516 3584
rect 2476 3516 2484 3524
rect 2492 3516 2500 3524
rect 2412 3496 2420 3504
rect 2412 3476 2420 3484
rect 2604 3796 2612 3804
rect 2700 4076 2708 4084
rect 2700 4056 2708 4064
rect 2652 3876 2660 3884
rect 2988 5056 2996 5064
rect 2988 4976 2996 4984
rect 3052 5296 3060 5304
rect 3180 5296 3188 5304
rect 3516 5336 3524 5344
rect 3308 5316 3316 5324
rect 3356 5316 3364 5324
rect 3420 5316 3428 5324
rect 3276 5296 3284 5304
rect 3404 5296 3412 5304
rect 3484 5296 3492 5304
rect 3292 5276 3300 5284
rect 3324 5276 3332 5284
rect 3500 5276 3508 5284
rect 3052 5136 3060 5144
rect 3148 5136 3156 5144
rect 3036 5096 3044 5104
rect 3420 5176 3428 5184
rect 3244 5136 3252 5144
rect 3260 5116 3268 5124
rect 3260 5096 3268 5104
rect 3020 5076 3028 5084
rect 3084 5076 3092 5084
rect 3164 5076 3172 5084
rect 3118 5006 3126 5014
rect 3132 5006 3140 5014
rect 3146 5006 3154 5014
rect 3052 4996 3060 5004
rect 3180 4996 3188 5004
rect 3116 4976 3124 4984
rect 3004 4956 3012 4964
rect 3052 4936 3060 4944
rect 2972 4916 2980 4924
rect 2972 4896 2980 4904
rect 3036 4896 3044 4904
rect 3052 4896 3060 4904
rect 3036 4836 3044 4844
rect 3020 4756 3028 4764
rect 3292 5016 3300 5024
rect 3324 5116 3332 5124
rect 3372 5116 3380 5124
rect 3404 5116 3412 5124
rect 3340 5076 3348 5084
rect 3324 5056 3332 5064
rect 3372 5056 3380 5064
rect 3388 5056 3396 5064
rect 3356 5016 3364 5024
rect 3372 4996 3380 5004
rect 3212 4976 3220 4984
rect 3276 4936 3284 4944
rect 3180 4856 3188 4864
rect 2908 4736 2916 4744
rect 2956 4736 2964 4744
rect 2988 4716 2996 4724
rect 2940 4696 2948 4704
rect 2956 4676 2964 4684
rect 2876 4596 2884 4604
rect 2860 4516 2868 4524
rect 2876 4396 2884 4404
rect 2812 4296 2820 4304
rect 2924 4536 2932 4544
rect 2972 4536 2980 4544
rect 2908 4476 2916 4484
rect 2892 4276 2900 4284
rect 2828 4196 2836 4204
rect 2860 4196 2868 4204
rect 2796 4176 2804 4184
rect 2812 4156 2820 4164
rect 2812 4096 2820 4104
rect 2780 4056 2788 4064
rect 2940 4496 2948 4504
rect 3020 4656 3028 4664
rect 2988 4496 2996 4504
rect 3020 4476 3028 4484
rect 3004 4456 3012 4464
rect 2956 4416 2964 4424
rect 3052 4736 3060 4744
rect 3084 4696 3092 4704
rect 3100 4676 3108 4684
rect 3052 4656 3060 4664
rect 3118 4606 3126 4614
rect 3132 4606 3140 4614
rect 3146 4606 3154 4614
rect 3180 4576 3188 4584
rect 3884 5736 3892 5744
rect 4060 5736 4068 5744
rect 4124 5736 4132 5744
rect 4140 5736 4148 5744
rect 4396 5756 4404 5764
rect 4444 5756 4452 5764
rect 4588 5756 4596 5764
rect 4220 5736 4228 5744
rect 4236 5736 4244 5744
rect 4444 5736 4452 5744
rect 4908 5776 4916 5784
rect 5004 5776 5012 5784
rect 5036 5776 5044 5784
rect 4988 5756 4996 5764
rect 4716 5736 4724 5744
rect 4092 5716 4100 5724
rect 4748 5716 4756 5724
rect 3596 5576 3604 5584
rect 3884 5576 3892 5584
rect 3772 5556 3780 5564
rect 3884 5556 3892 5564
rect 3628 5516 3636 5524
rect 3740 5516 3748 5524
rect 3676 5496 3684 5504
rect 3708 5496 3716 5504
rect 3580 5376 3588 5384
rect 3596 5376 3604 5384
rect 3868 5496 3876 5504
rect 4428 5696 4436 5704
rect 4508 5696 4516 5704
rect 4524 5696 4532 5704
rect 4604 5696 4612 5704
rect 4764 5696 4772 5704
rect 4844 5696 4852 5704
rect 4556 5676 4564 5684
rect 4732 5676 4740 5684
rect 4268 5656 4276 5664
rect 4284 5596 4292 5604
rect 4220 5536 4228 5544
rect 4252 5536 4260 5544
rect 4300 5536 4308 5544
rect 4380 5536 4388 5544
rect 4108 5516 4116 5524
rect 4284 5516 4292 5524
rect 3932 5496 3940 5504
rect 3692 5436 3700 5444
rect 3932 5476 3940 5484
rect 4044 5496 4052 5504
rect 4156 5496 4164 5504
rect 4316 5496 4324 5504
rect 3980 5476 3988 5484
rect 4060 5476 4068 5484
rect 3628 5316 3636 5324
rect 3532 5156 3540 5164
rect 3612 5156 3620 5164
rect 3436 5136 3444 5144
rect 3484 5136 3492 5144
rect 3532 5136 3540 5144
rect 3548 5136 3556 5144
rect 3452 5116 3460 5124
rect 3516 5096 3524 5104
rect 3500 5076 3508 5084
rect 3580 5096 3588 5104
rect 3564 5076 3572 5084
rect 3580 5076 3588 5084
rect 3420 5056 3428 5064
rect 3500 5036 3508 5044
rect 3564 5036 3572 5044
rect 3532 5016 3540 5024
rect 3452 4936 3460 4944
rect 3404 4916 3412 4924
rect 3468 4916 3476 4924
rect 3532 4916 3540 4924
rect 3388 4896 3396 4904
rect 3228 4876 3236 4884
rect 3404 4876 3412 4884
rect 3212 4856 3220 4864
rect 3228 4856 3236 4864
rect 3388 4836 3396 4844
rect 3372 4796 3380 4804
rect 3356 4736 3364 4744
rect 3260 4716 3268 4724
rect 3292 4716 3300 4724
rect 3340 4716 3348 4724
rect 3244 4696 3252 4704
rect 3228 4676 3236 4684
rect 3260 4676 3268 4684
rect 3212 4636 3220 4644
rect 3276 4636 3284 4644
rect 3228 4576 3236 4584
rect 3260 4576 3268 4584
rect 3068 4536 3076 4544
rect 3276 4536 3284 4544
rect 3052 4516 3060 4524
rect 3052 4496 3060 4504
rect 2988 4336 2996 4344
rect 2876 4076 2884 4084
rect 2748 3936 2756 3944
rect 2716 3916 2724 3924
rect 2780 3916 2788 3924
rect 2716 3896 2724 3904
rect 2764 3896 2772 3904
rect 2748 3876 2756 3884
rect 2668 3796 2676 3804
rect 2652 3736 2660 3744
rect 2588 3676 2596 3684
rect 2588 3596 2596 3604
rect 2556 3576 2564 3584
rect 2476 3476 2484 3484
rect 2492 3476 2500 3484
rect 2444 3456 2452 3464
rect 2460 3456 2468 3464
rect 2524 3396 2532 3404
rect 2444 3376 2452 3384
rect 2492 3376 2500 3384
rect 2508 3376 2516 3384
rect 2428 3356 2436 3364
rect 2492 3316 2500 3324
rect 2652 3616 2660 3624
rect 2620 3536 2628 3544
rect 2652 3536 2660 3544
rect 2716 3836 2724 3844
rect 2748 3836 2756 3844
rect 2780 3856 2788 3864
rect 2764 3816 2772 3824
rect 2764 3756 2772 3764
rect 2748 3716 2756 3724
rect 2732 3656 2740 3664
rect 2716 3556 2724 3564
rect 2588 3436 2596 3444
rect 2636 3396 2644 3404
rect 2572 3376 2580 3384
rect 2540 3356 2548 3364
rect 2556 3356 2564 3364
rect 2700 3516 2708 3524
rect 2684 3496 2692 3504
rect 2700 3456 2708 3464
rect 2748 3616 2756 3624
rect 2892 4036 2900 4044
rect 2844 3936 2852 3944
rect 2828 3916 2836 3924
rect 2812 3876 2820 3884
rect 2828 3836 2836 3844
rect 2844 3796 2852 3804
rect 2828 3776 2836 3784
rect 2812 3696 2820 3704
rect 2796 3636 2804 3644
rect 2764 3536 2772 3544
rect 2732 3516 2740 3524
rect 2780 3516 2788 3524
rect 2748 3496 2756 3504
rect 2780 3476 2788 3484
rect 2892 3836 2900 3844
rect 2892 3796 2900 3804
rect 2924 4196 2932 4204
rect 3004 4316 3012 4324
rect 2972 4196 2980 4204
rect 2956 4156 2964 4164
rect 2940 4116 2948 4124
rect 3164 4496 3172 4504
rect 3244 4496 3252 4504
rect 3148 4476 3156 4484
rect 3084 4436 3092 4444
rect 3180 4436 3188 4444
rect 3228 4436 3236 4444
rect 3068 4416 3076 4424
rect 3196 4396 3204 4404
rect 3308 4696 3316 4704
rect 3324 4676 3332 4684
rect 3324 4516 3332 4524
rect 3436 4896 3444 4904
rect 3516 4896 3524 4904
rect 3532 4896 3540 4904
rect 3500 4856 3508 4864
rect 3420 4836 3428 4844
rect 3468 4836 3476 4844
rect 3404 4796 3412 4804
rect 3500 4816 3508 4824
rect 3500 4736 3508 4744
rect 3420 4716 3428 4724
rect 3404 4696 3412 4704
rect 3436 4696 3444 4704
rect 3484 4676 3492 4684
rect 3548 4876 3556 4884
rect 3644 5116 3652 5124
rect 3628 5096 3636 5104
rect 3644 5076 3652 5084
rect 3660 5076 3668 5084
rect 3804 5436 3812 5444
rect 3948 5436 3956 5444
rect 3900 5416 3908 5424
rect 3740 5356 3748 5364
rect 3788 5336 3796 5344
rect 3740 5316 3748 5324
rect 3772 5316 3780 5324
rect 3884 5336 3892 5344
rect 3820 5316 3828 5324
rect 3868 5296 3876 5304
rect 3836 5276 3844 5284
rect 3804 5236 3812 5244
rect 3852 5236 3860 5244
rect 3932 5376 3940 5384
rect 3916 5196 3924 5204
rect 3948 5196 3956 5204
rect 3916 5176 3924 5184
rect 3740 5156 3748 5164
rect 3708 5136 3716 5144
rect 3868 5136 3876 5144
rect 3932 5136 3940 5144
rect 3708 5116 3716 5124
rect 3788 5116 3796 5124
rect 3692 5096 3700 5104
rect 3740 5096 3748 5104
rect 3724 5076 3732 5084
rect 3660 5056 3668 5064
rect 3676 5056 3684 5064
rect 3820 5076 3828 5084
rect 3788 5056 3796 5064
rect 3772 5036 3780 5044
rect 3804 4976 3812 4984
rect 3884 5116 3892 5124
rect 3852 5036 3860 5044
rect 3852 5016 3860 5024
rect 3900 5056 3908 5064
rect 3884 5036 3892 5044
rect 3820 4956 3828 4964
rect 3868 4956 3876 4964
rect 3916 4956 3924 4964
rect 3580 4916 3588 4924
rect 3996 5456 4004 5464
rect 4092 5436 4100 5444
rect 3996 5416 4004 5424
rect 3980 5336 3988 5344
rect 4124 5476 4132 5484
rect 4188 5480 4196 5484
rect 4188 5476 4196 5480
rect 4156 5456 4164 5464
rect 4268 5436 4276 5444
rect 4364 5476 4372 5484
rect 4380 5436 4388 5444
rect 4060 5376 4068 5384
rect 4316 5376 4324 5384
rect 4092 5356 4100 5364
rect 4140 5356 4148 5364
rect 4204 5356 4212 5364
rect 4284 5356 4292 5364
rect 4124 5316 4132 5324
rect 4300 5336 4308 5344
rect 4188 5316 4196 5324
rect 4220 5316 4228 5324
rect 4316 5316 4324 5324
rect 4108 5296 4116 5304
rect 4156 5296 4164 5304
rect 4284 5296 4292 5304
rect 4268 5176 4276 5184
rect 4638 5606 4646 5614
rect 4652 5606 4660 5614
rect 4666 5606 4674 5614
rect 4732 5576 4740 5584
rect 4604 5536 4612 5544
rect 4412 5516 4420 5524
rect 4476 5516 4484 5524
rect 4492 5516 4500 5524
rect 4604 5516 4612 5524
rect 4428 5476 4436 5484
rect 4460 5336 4468 5344
rect 4476 5316 4484 5324
rect 4572 5456 4580 5464
rect 4524 5436 4532 5444
rect 4508 5316 4516 5324
rect 4604 5456 4612 5464
rect 4636 5436 4644 5444
rect 4716 5496 4724 5504
rect 4748 5496 4756 5504
rect 4812 5676 4820 5684
rect 4796 5576 4804 5584
rect 4572 5316 4580 5324
rect 4924 5716 4932 5724
rect 4892 5696 4900 5704
rect 5148 5756 5156 5764
rect 5404 5756 5412 5764
rect 5452 5756 5460 5764
rect 5596 5756 5604 5764
rect 5164 5736 5172 5744
rect 5068 5716 5076 5724
rect 5116 5716 5124 5724
rect 4972 5696 4980 5704
rect 5020 5696 5028 5704
rect 5100 5676 5108 5684
rect 4956 5656 4964 5664
rect 5052 5656 5060 5664
rect 5036 5576 5044 5584
rect 4892 5536 4900 5544
rect 4940 5536 4948 5544
rect 4908 5516 4916 5524
rect 4908 5496 4916 5504
rect 4780 5436 4788 5444
rect 4844 5436 4852 5444
rect 4876 5436 4884 5444
rect 4956 5496 4964 5504
rect 5036 5496 5044 5504
rect 5020 5476 5028 5484
rect 4972 5456 4980 5464
rect 4924 5416 4932 5424
rect 4956 5416 4964 5424
rect 4988 5416 4996 5424
rect 5068 5496 5076 5504
rect 5132 5536 5140 5544
rect 5100 5496 5108 5504
rect 5084 5476 5092 5484
rect 4908 5376 4916 5384
rect 4972 5376 4980 5384
rect 4892 5356 4900 5364
rect 4924 5356 4932 5364
rect 4732 5336 4740 5344
rect 4892 5336 4900 5344
rect 4684 5316 4692 5324
rect 4796 5316 4804 5324
rect 4556 5296 4564 5304
rect 4700 5296 4708 5304
rect 4716 5256 4724 5264
rect 4460 5236 4468 5244
rect 4638 5206 4646 5214
rect 4652 5206 4660 5214
rect 4666 5206 4674 5214
rect 4908 5316 4916 5324
rect 4972 5316 4980 5324
rect 5036 5316 5044 5324
rect 4860 5296 4868 5304
rect 4892 5296 4900 5304
rect 4492 5176 4500 5184
rect 4524 5176 4532 5184
rect 4188 5156 4196 5164
rect 4396 5156 4404 5164
rect 4476 5156 4484 5164
rect 4076 5116 4084 5124
rect 4140 5116 4148 5124
rect 3964 5096 3972 5104
rect 4060 5096 4068 5104
rect 3980 5076 3988 5084
rect 4044 5076 4052 5084
rect 3964 5036 3972 5044
rect 3980 5036 3988 5044
rect 3788 4916 3796 4924
rect 3836 4916 3844 4924
rect 3612 4896 3620 4904
rect 3644 4896 3652 4904
rect 3596 4876 3604 4884
rect 3644 4876 3652 4884
rect 3564 4736 3572 4744
rect 3708 4876 3716 4884
rect 3676 4856 3684 4864
rect 3740 4856 3748 4864
rect 3660 4836 3668 4844
rect 3724 4836 3732 4844
rect 3772 4816 3780 4824
rect 3852 4816 3860 4824
rect 3900 4916 3908 4924
rect 3996 5016 4004 5024
rect 3996 4956 4004 4964
rect 3980 4936 3988 4944
rect 3948 4916 3956 4924
rect 3964 4896 3972 4904
rect 3644 4776 3652 4784
rect 3788 4776 3796 4784
rect 3884 4776 3892 4784
rect 3772 4756 3780 4764
rect 3756 4736 3764 4744
rect 3404 4656 3412 4664
rect 3452 4656 3460 4664
rect 3436 4636 3444 4644
rect 3404 4616 3412 4624
rect 3372 4496 3380 4504
rect 3388 4496 3396 4504
rect 3308 4476 3316 4484
rect 3340 4476 3348 4484
rect 3308 4456 3316 4464
rect 3180 4376 3188 4384
rect 3260 4376 3268 4384
rect 3164 4356 3172 4364
rect 3052 4316 3060 4324
rect 3036 4276 3044 4284
rect 3164 4316 3172 4324
rect 3180 4296 3188 4304
rect 3356 4416 3364 4424
rect 3468 4516 3476 4524
rect 3500 4516 3508 4524
rect 3420 4496 3428 4504
rect 3452 4496 3460 4504
rect 3436 4416 3444 4424
rect 3356 4356 3364 4364
rect 3340 4336 3348 4344
rect 3228 4316 3236 4324
rect 3148 4276 3156 4284
rect 3212 4276 3220 4284
rect 3260 4296 3268 4304
rect 3244 4236 3252 4244
rect 3118 4206 3126 4214
rect 3132 4206 3140 4214
rect 3146 4206 3154 4214
rect 3132 4176 3140 4184
rect 3084 4136 3092 4144
rect 2940 4096 2948 4104
rect 3004 4096 3012 4104
rect 2924 4016 2932 4024
rect 2924 3836 2932 3844
rect 2908 3776 2916 3784
rect 2988 4056 2996 4064
rect 2972 4036 2980 4044
rect 2956 3916 2964 3924
rect 2972 3896 2980 3904
rect 2956 3776 2964 3784
rect 2924 3736 2932 3744
rect 2924 3696 2932 3704
rect 2876 3636 2884 3644
rect 2924 3596 2932 3604
rect 2972 3736 2980 3744
rect 3004 3876 3012 3884
rect 3004 3736 3012 3744
rect 3052 4056 3060 4064
rect 3100 4076 3108 4084
rect 3068 4036 3076 4044
rect 3052 3916 3060 3924
rect 3068 3916 3076 3924
rect 3228 4136 3236 4144
rect 3196 4116 3204 4124
rect 3180 4096 3188 4104
rect 3244 4096 3252 4104
rect 3276 4176 3284 4184
rect 3276 4156 3284 4164
rect 3164 4036 3172 4044
rect 3276 4076 3284 4084
rect 3468 4436 3476 4444
rect 3516 4476 3524 4484
rect 3500 4456 3508 4464
rect 3388 4336 3396 4344
rect 3452 4336 3460 4344
rect 3308 4196 3316 4204
rect 3308 4136 3316 4144
rect 3420 4316 3428 4324
rect 3388 4296 3396 4304
rect 3436 4296 3444 4304
rect 3404 4276 3412 4284
rect 3452 4276 3460 4284
rect 3420 4236 3428 4244
rect 3356 4156 3364 4164
rect 3500 4316 3508 4324
rect 3484 4296 3492 4304
rect 3516 4256 3524 4264
rect 3548 4676 3556 4684
rect 3548 4656 3556 4664
rect 3836 4736 3844 4744
rect 3772 4716 3780 4724
rect 3820 4716 3828 4724
rect 3852 4716 3860 4724
rect 3884 4716 3892 4724
rect 3724 4696 3732 4704
rect 3756 4696 3764 4704
rect 3788 4696 3796 4704
rect 3660 4656 3668 4664
rect 3740 4676 3748 4684
rect 3644 4616 3652 4624
rect 3676 4616 3684 4624
rect 3724 4656 3732 4664
rect 3564 4596 3572 4604
rect 3628 4596 3636 4604
rect 3692 4596 3700 4604
rect 3548 4416 3556 4424
rect 3772 4656 3780 4664
rect 3612 4576 3620 4584
rect 3756 4576 3764 4584
rect 3836 4696 3844 4704
rect 3948 4696 3956 4704
rect 3932 4676 3940 4684
rect 3836 4656 3844 4664
rect 3900 4636 3908 4644
rect 3932 4616 3940 4624
rect 4028 4916 4036 4924
rect 4076 4976 4084 4984
rect 4060 4936 4068 4944
rect 4092 4956 4100 4964
rect 4156 5096 4164 5104
rect 4172 5076 4180 5084
rect 4300 5136 4308 5144
rect 4204 5116 4212 5124
rect 4236 5096 4244 5104
rect 4220 5076 4228 5084
rect 4700 5136 4708 5144
rect 4748 5136 4756 5144
rect 4828 5136 4836 5144
rect 4300 5116 4308 5124
rect 4332 5116 4340 5124
rect 4428 5116 4436 5124
rect 4460 5116 4468 5124
rect 4540 5116 4548 5124
rect 4300 5096 4308 5104
rect 4364 5096 4372 5104
rect 4284 5076 4292 5084
rect 4348 5076 4356 5084
rect 4380 5076 4388 5084
rect 4204 5056 4212 5064
rect 4252 5056 4260 5064
rect 4284 5056 4292 5064
rect 4236 5036 4244 5044
rect 4220 5016 4228 5024
rect 4140 4956 4148 4964
rect 4092 4916 4100 4924
rect 4140 4916 4148 4924
rect 4476 5096 4484 5104
rect 4540 5096 4548 5104
rect 4396 5056 4404 5064
rect 4428 5056 4436 5064
rect 4348 5036 4356 5044
rect 4268 4956 4276 4964
rect 4300 4956 4308 4964
rect 4364 4956 4372 4964
rect 4428 4956 4436 4964
rect 4204 4916 4212 4924
rect 4252 4916 4260 4924
rect 4332 4936 4340 4944
rect 4412 4936 4420 4944
rect 4316 4916 4324 4924
rect 4396 4916 4404 4924
rect 4044 4896 4052 4904
rect 4012 4776 4020 4784
rect 4076 4756 4084 4764
rect 4060 4736 4068 4744
rect 4012 4716 4020 4724
rect 4012 4696 4020 4704
rect 4140 4716 4148 4724
rect 4060 4696 4068 4704
rect 4108 4696 4116 4704
rect 4124 4696 4132 4704
rect 4108 4616 4116 4624
rect 4044 4596 4052 4604
rect 3852 4576 3860 4584
rect 4060 4576 4068 4584
rect 4140 4576 4148 4584
rect 3868 4556 3876 4564
rect 4012 4556 4020 4564
rect 3644 4536 3652 4544
rect 3884 4536 3892 4544
rect 3932 4536 3940 4544
rect 3980 4536 3988 4544
rect 3580 4516 3588 4524
rect 3612 4516 3620 4524
rect 3596 4496 3604 4504
rect 3628 4476 3636 4484
rect 3596 4456 3604 4464
rect 3580 4376 3588 4384
rect 3532 4236 3540 4244
rect 3532 4216 3540 4224
rect 3580 4256 3588 4264
rect 3564 4196 3572 4204
rect 3500 4176 3508 4184
rect 3548 4176 3556 4184
rect 3564 4176 3572 4184
rect 3372 4136 3380 4144
rect 3388 4136 3396 4144
rect 3436 4136 3444 4144
rect 3340 4096 3348 4104
rect 3404 4056 3412 4064
rect 3324 4016 3332 4024
rect 3420 4016 3428 4024
rect 3340 3976 3348 3984
rect 3420 3956 3428 3964
rect 3388 3936 3396 3944
rect 3404 3936 3412 3944
rect 3468 3936 3476 3944
rect 3484 3936 3492 3944
rect 3148 3916 3156 3924
rect 3196 3916 3204 3924
rect 3276 3916 3284 3924
rect 3036 3896 3044 3904
rect 3180 3896 3188 3904
rect 3244 3896 3252 3904
rect 3004 3676 3012 3684
rect 3004 3616 3012 3624
rect 2972 3576 2980 3584
rect 2924 3536 2932 3544
rect 2940 3536 2948 3544
rect 2988 3556 2996 3564
rect 3084 3816 3092 3824
rect 3052 3796 3060 3804
rect 3052 3756 3060 3764
rect 3118 3806 3126 3814
rect 3132 3806 3140 3814
rect 3146 3806 3154 3814
rect 3084 3736 3092 3744
rect 3068 3716 3076 3724
rect 3084 3696 3092 3704
rect 3084 3676 3092 3684
rect 3036 3616 3044 3624
rect 3036 3556 3044 3564
rect 3052 3556 3060 3564
rect 3020 3516 3028 3524
rect 3212 3856 3220 3864
rect 3340 3896 3348 3904
rect 3308 3876 3316 3884
rect 3324 3876 3332 3884
rect 3196 3816 3204 3824
rect 3244 3816 3252 3824
rect 3276 3816 3284 3824
rect 3356 3816 3364 3824
rect 3372 3816 3380 3824
rect 3324 3776 3332 3784
rect 3340 3776 3348 3784
rect 3180 3736 3188 3744
rect 3212 3716 3220 3724
rect 3116 3676 3124 3684
rect 3116 3636 3124 3644
rect 2972 3496 2980 3504
rect 3020 3496 3028 3504
rect 2940 3476 2948 3484
rect 3004 3476 3012 3484
rect 2716 3336 2724 3344
rect 2540 3316 2548 3324
rect 2620 3316 2628 3324
rect 2652 3316 2660 3324
rect 2444 3296 2452 3304
rect 2492 3296 2500 3304
rect 2428 3276 2436 3284
rect 2476 3276 2484 3284
rect 2636 3296 2644 3304
rect 2668 3296 2676 3304
rect 2524 3276 2532 3284
rect 2604 3276 2612 3284
rect 2412 3196 2420 3204
rect 2556 3176 2564 3184
rect 2396 3096 2404 3104
rect 2284 3056 2292 3064
rect 2156 2976 2164 2984
rect 2188 2956 2196 2964
rect 2380 3056 2388 3064
rect 2460 3096 2468 3104
rect 2444 3076 2452 3084
rect 2540 3076 2548 3084
rect 2316 3036 2324 3044
rect 2316 3016 2324 3024
rect 2300 2976 2308 2984
rect 2124 2936 2132 2944
rect 2284 2936 2292 2944
rect 2108 2916 2116 2924
rect 2268 2916 2276 2924
rect 2108 2896 2116 2904
rect 2044 2856 2052 2864
rect 1900 2836 1908 2844
rect 1948 2836 1956 2844
rect 1756 2776 1764 2784
rect 1676 2696 1684 2704
rect 1708 2696 1716 2704
rect 1740 2696 1748 2704
rect 1660 2676 1668 2684
rect 1692 2676 1700 2684
rect 1788 2736 1796 2744
rect 1996 2736 2004 2744
rect 1884 2716 1892 2724
rect 2028 2716 2036 2724
rect 1852 2696 1860 2704
rect 1772 2636 1780 2644
rect 1740 2616 1748 2624
rect 1580 2576 1588 2584
rect 1900 2696 1908 2704
rect 1964 2696 1972 2704
rect 1884 2676 1892 2684
rect 1980 2676 1988 2684
rect 1820 2636 1828 2644
rect 1948 2636 1956 2644
rect 1804 2576 1812 2584
rect 1660 2536 1668 2544
rect 1708 2536 1716 2544
rect 1788 2536 1796 2544
rect 1612 2516 1620 2524
rect 1692 2516 1700 2524
rect 1516 2476 1524 2484
rect 1500 2296 1508 2304
rect 1884 2596 1892 2604
rect 1996 2596 2004 2604
rect 1868 2576 1876 2584
rect 1740 2516 1748 2524
rect 1916 2556 1924 2564
rect 1948 2556 1956 2564
rect 1580 2496 1588 2504
rect 1900 2496 1908 2504
rect 1548 2476 1556 2484
rect 1692 2476 1700 2484
rect 1566 2406 1574 2414
rect 1580 2406 1588 2414
rect 1594 2406 1602 2414
rect 1644 2396 1652 2404
rect 1532 2296 1540 2304
rect 1564 2296 1572 2304
rect 1516 2276 1524 2284
rect 1676 2336 1684 2344
rect 1372 2236 1380 2244
rect 1420 2236 1428 2244
rect 1356 2216 1364 2224
rect 1340 2136 1348 2144
rect 1660 2256 1668 2264
rect 1500 2196 1508 2204
rect 1532 2216 1540 2224
rect 1404 2176 1412 2184
rect 1436 2176 1444 2184
rect 1516 2176 1524 2184
rect 1516 2156 1524 2164
rect 1276 2096 1284 2104
rect 1308 2096 1316 2104
rect 1260 2076 1268 2084
rect 1404 2136 1412 2144
rect 1420 2116 1428 2124
rect 1500 2116 1508 2124
rect 1676 2156 1684 2164
rect 1628 2116 1636 2124
rect 1644 2116 1652 2124
rect 1660 2116 1668 2124
rect 1324 2076 1332 2084
rect 1292 2036 1300 2044
rect 1276 1996 1284 2004
rect 1356 1976 1364 1984
rect 1340 1956 1348 1964
rect 1260 1936 1268 1944
rect 1324 1936 1332 1944
rect 1292 1896 1300 1904
rect 1324 1896 1332 1904
rect 1276 1856 1284 1864
rect 1180 1716 1188 1724
rect 1116 1656 1124 1664
rect 1132 1656 1140 1664
rect 1148 1636 1156 1644
rect 1100 1556 1108 1564
rect 1084 1536 1092 1544
rect 1100 1536 1108 1544
rect 1020 1496 1028 1504
rect 1068 1496 1076 1504
rect 1100 1496 1108 1504
rect 988 1476 996 1484
rect 1084 1476 1092 1484
rect 1068 1456 1076 1464
rect 1020 1436 1028 1444
rect 1052 1416 1060 1424
rect 972 1396 980 1404
rect 1020 1396 1028 1404
rect 956 1376 964 1384
rect 956 1356 964 1364
rect 1180 1596 1188 1604
rect 1196 1596 1204 1604
rect 1164 1556 1172 1564
rect 1196 1536 1204 1544
rect 1132 1476 1140 1484
rect 1100 1376 1108 1384
rect 972 1316 980 1324
rect 988 1316 996 1324
rect 892 1296 900 1304
rect 940 1296 948 1304
rect 956 1296 964 1304
rect 1020 1296 1028 1304
rect 1052 1296 1060 1304
rect 876 1276 884 1284
rect 860 1156 868 1164
rect 812 1116 820 1124
rect 844 1096 852 1104
rect 764 976 772 984
rect 732 956 740 964
rect 860 1056 868 1064
rect 924 1236 932 1244
rect 908 1196 916 1204
rect 988 1216 996 1224
rect 940 1176 948 1184
rect 972 1176 980 1184
rect 1164 1456 1172 1464
rect 1148 1396 1156 1404
rect 1132 1256 1140 1264
rect 1084 1216 1092 1224
rect 1004 1156 1012 1164
rect 1068 1156 1076 1164
rect 908 1076 916 1084
rect 956 1076 964 1084
rect 972 1076 980 1084
rect 988 1056 996 1064
rect 796 976 804 984
rect 844 976 852 984
rect 812 956 820 964
rect 748 936 756 944
rect 780 936 788 944
rect 636 916 644 924
rect 652 916 660 924
rect 620 896 628 904
rect 252 876 260 884
rect 396 876 404 884
rect 556 876 564 884
rect 604 876 612 884
rect 620 836 628 844
rect 236 776 244 784
rect 252 716 260 724
rect 300 776 308 784
rect 332 776 340 784
rect 172 696 180 704
rect 204 696 212 704
rect 284 696 292 704
rect 204 676 212 684
rect 220 676 228 684
rect 108 616 116 624
rect 92 576 100 584
rect 92 556 100 564
rect 108 536 116 544
rect 220 616 228 624
rect 140 576 148 584
rect 204 576 212 584
rect 252 596 260 604
rect 316 756 324 764
rect 316 736 324 744
rect 364 736 372 744
rect 492 776 500 784
rect 588 776 596 784
rect 380 716 388 724
rect 412 736 420 744
rect 428 736 436 744
rect 460 736 468 744
rect 492 736 500 744
rect 540 736 548 744
rect 348 696 356 704
rect 428 696 436 704
rect 364 656 372 664
rect 396 656 404 664
rect 332 576 340 584
rect 380 536 388 544
rect 268 516 276 524
rect 316 516 324 524
rect 188 496 196 504
rect 236 496 244 504
rect 332 496 340 504
rect 140 476 148 484
rect 284 476 292 484
rect 300 476 308 484
rect 236 456 244 464
rect 76 436 84 444
rect 124 436 132 444
rect 44 376 52 384
rect 124 416 132 424
rect 92 376 100 384
rect 44 316 52 324
rect 60 296 68 304
rect 140 316 148 324
rect 204 316 212 324
rect 412 476 420 484
rect 396 416 404 424
rect 300 396 308 404
rect 348 396 356 404
rect 396 396 404 404
rect 268 356 276 364
rect 252 336 260 344
rect 124 296 132 304
rect 156 296 164 304
rect 220 296 228 304
rect 44 276 52 284
rect 92 276 100 284
rect 204 276 212 284
rect 188 256 196 264
rect 76 156 84 164
rect 172 216 180 224
rect 140 196 148 204
rect 252 276 260 284
rect 316 296 324 304
rect 364 296 372 304
rect 380 276 388 284
rect 412 276 420 284
rect 236 256 244 264
rect 364 256 372 264
rect 524 696 532 704
rect 572 696 580 704
rect 668 856 676 864
rect 652 756 660 764
rect 620 696 628 704
rect 444 676 452 684
rect 508 676 516 684
rect 588 656 596 664
rect 636 656 644 664
rect 524 596 532 604
rect 620 596 628 604
rect 604 576 612 584
rect 460 556 468 564
rect 508 556 516 564
rect 572 556 580 564
rect 492 496 500 504
rect 572 516 580 524
rect 540 496 548 504
rect 652 636 660 644
rect 684 836 692 844
rect 684 716 692 724
rect 828 736 836 744
rect 780 696 788 704
rect 828 696 836 704
rect 764 676 772 684
rect 812 676 820 684
rect 844 676 852 684
rect 684 596 692 604
rect 780 656 788 664
rect 796 616 804 624
rect 684 576 692 584
rect 716 576 724 584
rect 732 576 740 584
rect 764 576 772 584
rect 780 576 788 584
rect 636 556 644 564
rect 700 556 708 564
rect 636 536 644 544
rect 700 536 708 544
rect 732 536 740 544
rect 748 516 756 524
rect 476 476 484 484
rect 524 476 532 484
rect 684 476 692 484
rect 716 476 724 484
rect 732 476 740 484
rect 780 476 788 484
rect 444 436 452 444
rect 492 416 500 424
rect 460 376 468 384
rect 444 296 452 304
rect 348 236 356 244
rect 236 216 244 224
rect 220 176 228 184
rect 188 136 196 144
rect 76 116 84 124
rect 188 116 196 124
rect 44 98 52 104
rect 44 96 52 98
rect 540 396 548 404
rect 556 356 564 364
rect 492 336 500 344
rect 588 336 596 344
rect 476 316 484 324
rect 508 296 516 304
rect 572 316 580 324
rect 556 296 564 304
rect 684 396 692 404
rect 700 396 708 404
rect 636 316 644 324
rect 652 316 660 324
rect 620 296 628 304
rect 684 296 692 304
rect 652 256 660 264
rect 428 216 436 224
rect 412 196 420 204
rect 540 236 548 244
rect 604 236 612 244
rect 460 196 468 204
rect 524 176 532 184
rect 588 176 596 184
rect 284 156 292 164
rect 252 116 260 124
rect 316 116 324 124
rect 364 136 372 144
rect 380 136 388 144
rect 540 156 548 164
rect 508 136 516 144
rect 556 136 564 144
rect 396 116 404 124
rect 444 116 452 124
rect 492 116 500 124
rect 668 196 676 204
rect 828 596 836 604
rect 940 1036 948 1044
rect 892 1016 900 1024
rect 972 1016 980 1024
rect 908 996 916 1004
rect 940 956 948 964
rect 908 876 916 884
rect 924 796 932 804
rect 988 876 996 884
rect 940 756 948 764
rect 972 756 980 764
rect 940 716 948 724
rect 924 676 932 684
rect 988 676 996 684
rect 1068 1116 1076 1124
rect 1052 1096 1060 1104
rect 1052 1056 1060 1064
rect 1036 1036 1044 1044
rect 1020 1016 1028 1024
rect 1020 996 1028 1004
rect 1036 976 1044 984
rect 1068 956 1076 964
rect 1116 1136 1124 1144
rect 1116 1036 1124 1044
rect 1084 916 1092 924
rect 1212 1456 1220 1464
rect 1244 1736 1252 1744
rect 1308 1736 1316 1744
rect 1372 1936 1380 1944
rect 1356 1916 1364 1924
rect 1372 1916 1380 1924
rect 1356 1876 1364 1884
rect 1628 2096 1636 2104
rect 1644 2076 1652 2084
rect 1420 2056 1428 2064
rect 1500 2056 1508 2064
rect 1452 2016 1460 2024
rect 1660 2016 1668 2024
rect 1436 1976 1444 1984
rect 1420 1936 1428 1944
rect 1388 1856 1396 1864
rect 1404 1836 1412 1844
rect 1566 2006 1574 2014
rect 1580 2006 1588 2014
rect 1594 2006 1602 2014
rect 1644 1996 1652 2004
rect 1564 1956 1572 1964
rect 1452 1916 1460 1924
rect 1500 1916 1508 1924
rect 1516 1896 1524 1904
rect 1436 1876 1444 1884
rect 1484 1876 1492 1884
rect 1420 1796 1428 1804
rect 1372 1776 1380 1784
rect 1420 1776 1428 1784
rect 1244 1716 1252 1724
rect 1292 1716 1300 1724
rect 1340 1716 1348 1724
rect 1644 1856 1652 1864
rect 1516 1816 1524 1824
rect 1452 1796 1460 1804
rect 1468 1796 1476 1804
rect 1356 1696 1364 1704
rect 1372 1696 1380 1704
rect 1260 1656 1268 1664
rect 1324 1656 1332 1664
rect 1356 1656 1364 1664
rect 1276 1596 1284 1604
rect 1260 1576 1268 1584
rect 1244 1496 1252 1504
rect 1292 1556 1300 1564
rect 1292 1536 1300 1544
rect 1308 1496 1316 1504
rect 1228 1396 1236 1404
rect 1212 1376 1220 1384
rect 1196 1336 1204 1344
rect 1244 1336 1252 1344
rect 1212 1316 1220 1324
rect 1228 1316 1236 1324
rect 1244 1296 1252 1304
rect 1180 1276 1188 1284
rect 1180 1136 1188 1144
rect 1164 1076 1172 1084
rect 1148 976 1156 984
rect 1148 916 1156 924
rect 1068 896 1076 904
rect 1100 896 1108 904
rect 1132 896 1140 904
rect 1020 876 1028 884
rect 1084 876 1092 884
rect 1276 1436 1284 1444
rect 1292 1376 1300 1384
rect 1276 1336 1284 1344
rect 1260 1176 1268 1184
rect 1228 1136 1236 1144
rect 1212 996 1220 1004
rect 1196 916 1204 924
rect 1116 876 1124 884
rect 1164 876 1172 884
rect 1100 816 1108 824
rect 1100 796 1108 804
rect 1020 776 1028 784
rect 1036 736 1044 744
rect 1148 796 1156 804
rect 1116 776 1124 784
rect 1132 776 1140 784
rect 1068 716 1076 724
rect 1180 816 1188 824
rect 1164 716 1172 724
rect 1068 676 1076 684
rect 1164 676 1172 684
rect 1340 1576 1348 1584
rect 1388 1636 1396 1644
rect 1356 1496 1364 1504
rect 1372 1456 1380 1464
rect 1356 1396 1364 1404
rect 1356 1376 1364 1384
rect 1628 1796 1636 1804
rect 1548 1776 1556 1784
rect 1484 1736 1492 1744
rect 1500 1736 1508 1744
rect 1532 1736 1540 1744
rect 1468 1716 1476 1724
rect 1468 1676 1476 1684
rect 1452 1556 1460 1564
rect 1596 1736 1604 1744
rect 1548 1676 1556 1684
rect 1612 1656 1620 1664
rect 1532 1636 1540 1644
rect 1516 1616 1524 1624
rect 1566 1606 1574 1614
rect 1580 1606 1588 1614
rect 1594 1606 1602 1614
rect 1532 1596 1540 1604
rect 1500 1576 1508 1584
rect 1564 1556 1572 1564
rect 1500 1536 1508 1544
rect 1548 1516 1556 1524
rect 1484 1496 1492 1504
rect 1404 1416 1412 1424
rect 1436 1416 1444 1424
rect 1420 1396 1428 1404
rect 1468 1376 1476 1384
rect 1340 1336 1348 1344
rect 1452 1336 1460 1344
rect 1580 1456 1588 1464
rect 1580 1356 1588 1364
rect 1724 2376 1732 2384
rect 1836 2376 1844 2384
rect 1724 2356 1732 2364
rect 1772 2356 1780 2364
rect 1852 2356 1860 2364
rect 1740 2316 1748 2324
rect 1804 2336 1812 2344
rect 1836 2336 1844 2344
rect 1708 2276 1716 2284
rect 1788 2276 1796 2284
rect 1820 2316 1828 2324
rect 2092 2736 2100 2744
rect 2172 2876 2180 2884
rect 2140 2856 2148 2864
rect 2172 2756 2180 2764
rect 2268 2896 2276 2904
rect 2300 2856 2308 2864
rect 2284 2756 2292 2764
rect 2188 2736 2196 2744
rect 2220 2736 2228 2744
rect 2076 2696 2084 2704
rect 2108 2696 2116 2704
rect 2060 2676 2068 2684
rect 2172 2696 2180 2704
rect 2204 2696 2212 2704
rect 2332 2916 2340 2924
rect 2348 2896 2356 2904
rect 2412 2916 2420 2924
rect 2396 2896 2404 2904
rect 2380 2876 2388 2884
rect 2428 2876 2436 2884
rect 2332 2756 2340 2764
rect 2380 2756 2388 2764
rect 2284 2696 2292 2704
rect 2252 2676 2260 2684
rect 2300 2676 2308 2684
rect 2476 3016 2484 3024
rect 2508 3016 2516 3024
rect 2700 3296 2708 3304
rect 2684 3256 2692 3264
rect 2716 3256 2724 3264
rect 2604 3176 2612 3184
rect 2604 3156 2612 3164
rect 2636 3156 2644 3164
rect 2796 3456 2804 3464
rect 2892 3436 2900 3444
rect 2940 3436 2948 3444
rect 2988 3436 2996 3444
rect 2764 3396 2772 3404
rect 2828 3396 2836 3404
rect 2748 3356 2756 3364
rect 2812 3356 2820 3364
rect 2796 3336 2804 3344
rect 2860 3376 2868 3384
rect 2844 3356 2852 3364
rect 2876 3336 2884 3344
rect 2908 3336 2916 3344
rect 2844 3316 2852 3324
rect 2780 3276 2788 3284
rect 2812 3276 2820 3284
rect 2700 3176 2708 3184
rect 2684 3136 2692 3144
rect 2588 3096 2596 3104
rect 2652 3096 2660 3104
rect 2668 3076 2676 3084
rect 2572 2996 2580 3004
rect 2620 2996 2628 3004
rect 2588 2976 2596 2984
rect 2508 2956 2516 2964
rect 2572 2956 2580 2964
rect 2540 2916 2548 2924
rect 2492 2896 2500 2904
rect 2748 3156 2756 3164
rect 2812 3136 2820 3144
rect 2764 3116 2772 3124
rect 2684 2976 2692 2984
rect 2652 2956 2660 2964
rect 2700 2916 2708 2924
rect 2860 3176 2868 3184
rect 2924 3316 2932 3324
rect 2924 3216 2932 3224
rect 2908 3156 2916 3164
rect 2860 3136 2868 3144
rect 2892 3136 2900 3144
rect 2844 3116 2852 3124
rect 2828 3096 2836 3104
rect 2876 3096 2884 3104
rect 2748 3076 2756 3084
rect 2876 3076 2884 3084
rect 2844 3056 2852 3064
rect 2812 3036 2820 3044
rect 2796 2956 2804 2964
rect 2732 2936 2740 2944
rect 2732 2916 2740 2924
rect 2748 2916 2756 2924
rect 2460 2876 2468 2884
rect 2524 2876 2532 2884
rect 2444 2816 2452 2824
rect 2412 2736 2420 2744
rect 2460 2736 2468 2744
rect 2428 2716 2436 2724
rect 2428 2696 2436 2704
rect 2348 2676 2356 2684
rect 2668 2876 2676 2884
rect 2620 2836 2628 2844
rect 2636 2816 2644 2824
rect 2588 2716 2596 2724
rect 2620 2716 2628 2724
rect 2476 2696 2484 2704
rect 2604 2696 2612 2704
rect 2476 2676 2484 2684
rect 2060 2656 2068 2664
rect 2172 2656 2180 2664
rect 2236 2656 2244 2664
rect 2316 2656 2324 2664
rect 2380 2656 2388 2664
rect 2444 2656 2452 2664
rect 2492 2656 2500 2664
rect 2108 2576 2116 2584
rect 2012 2556 2020 2564
rect 2012 2536 2020 2544
rect 2124 2556 2132 2564
rect 1980 2496 1988 2504
rect 2076 2496 2084 2504
rect 1996 2476 2004 2484
rect 1964 2456 1972 2464
rect 1948 2396 1956 2404
rect 1900 2356 1908 2364
rect 2124 2456 2132 2464
rect 2060 2396 2068 2404
rect 1996 2376 2004 2384
rect 1980 2356 1988 2364
rect 1900 2336 1908 2344
rect 1884 2316 1892 2324
rect 1932 2316 1940 2324
rect 1948 2316 1956 2324
rect 1884 2276 1892 2284
rect 1868 2216 1876 2224
rect 1724 2196 1732 2204
rect 1708 2116 1716 2124
rect 2092 2376 2100 2384
rect 2012 2316 2020 2324
rect 2044 2316 2052 2324
rect 2156 2536 2164 2544
rect 2268 2636 2276 2644
rect 2236 2616 2244 2624
rect 2396 2616 2404 2624
rect 2300 2576 2308 2584
rect 2364 2576 2372 2584
rect 2316 2556 2324 2564
rect 2268 2516 2276 2524
rect 2220 2496 2228 2504
rect 2140 2336 2148 2344
rect 2188 2456 2196 2464
rect 2172 2396 2180 2404
rect 2380 2536 2388 2544
rect 2412 2536 2420 2544
rect 2428 2516 2436 2524
rect 2444 2516 2452 2524
rect 2332 2456 2340 2464
rect 2524 2636 2532 2644
rect 2588 2636 2596 2644
rect 2620 2616 2628 2624
rect 2652 2776 2660 2784
rect 2828 2896 2836 2904
rect 2748 2876 2756 2884
rect 2764 2876 2772 2884
rect 2748 2856 2756 2864
rect 2716 2816 2724 2824
rect 2732 2756 2740 2764
rect 2748 2756 2756 2764
rect 2668 2716 2676 2724
rect 2700 2716 2708 2724
rect 2700 2696 2708 2704
rect 2684 2656 2692 2664
rect 2652 2636 2660 2644
rect 2684 2636 2692 2644
rect 2524 2536 2532 2544
rect 2668 2536 2676 2544
rect 2508 2516 2516 2524
rect 2572 2516 2580 2524
rect 2652 2516 2660 2524
rect 2476 2496 2484 2504
rect 2492 2496 2500 2504
rect 2668 2496 2676 2504
rect 2460 2476 2468 2484
rect 2252 2436 2260 2444
rect 2348 2436 2356 2444
rect 2364 2436 2372 2444
rect 2268 2416 2276 2424
rect 2348 2396 2356 2404
rect 2268 2376 2276 2384
rect 2204 2356 2212 2364
rect 2316 2336 2324 2344
rect 1932 2256 1940 2264
rect 2108 2256 2116 2264
rect 1948 2236 1956 2244
rect 1996 2196 2004 2204
rect 2012 2156 2020 2164
rect 2028 2156 2036 2164
rect 1820 2136 1828 2144
rect 1884 2136 1892 2144
rect 1900 2136 1908 2144
rect 1964 2136 1972 2144
rect 1756 2096 1764 2104
rect 1852 2096 1860 2104
rect 1900 2096 1908 2104
rect 2092 2156 2100 2164
rect 2140 2176 2148 2184
rect 2172 2176 2180 2184
rect 2060 2136 2068 2144
rect 2012 2116 2020 2124
rect 2044 2116 2052 2124
rect 1948 2096 1956 2104
rect 1996 2096 2004 2104
rect 2028 2096 2036 2104
rect 2204 2276 2212 2284
rect 2476 2376 2484 2384
rect 2396 2336 2404 2344
rect 2460 2336 2468 2344
rect 2412 2316 2420 2324
rect 2476 2316 2484 2324
rect 2268 2296 2276 2304
rect 2252 2276 2260 2284
rect 2316 2276 2324 2284
rect 2364 2276 2372 2284
rect 2412 2276 2420 2284
rect 2236 2236 2244 2244
rect 2252 2236 2260 2244
rect 2428 2256 2436 2264
rect 2412 2216 2420 2224
rect 2316 2196 2324 2204
rect 2188 2156 2196 2164
rect 2300 2156 2308 2164
rect 2124 2116 2132 2124
rect 2156 2116 2164 2124
rect 2076 2096 2084 2104
rect 2204 2116 2212 2124
rect 2268 2116 2276 2124
rect 2252 2096 2260 2104
rect 1804 2076 1812 2084
rect 1868 2076 1876 2084
rect 1916 2076 1924 2084
rect 2252 2076 2260 2084
rect 1724 2056 1732 2064
rect 1900 2056 1908 2064
rect 2236 2056 2244 2064
rect 2300 2056 2308 2064
rect 1692 2016 1700 2024
rect 1676 1956 1684 1964
rect 1756 1976 1764 1984
rect 1724 1956 1732 1964
rect 1724 1916 1732 1924
rect 1740 1896 1748 1904
rect 1692 1876 1700 1884
rect 1724 1876 1732 1884
rect 1756 1876 1764 1884
rect 1868 1996 1876 2004
rect 2012 2036 2020 2044
rect 1948 1996 1956 2004
rect 1804 1916 1812 1924
rect 1868 1916 1876 1924
rect 1900 1916 1908 1924
rect 1932 1916 1940 1924
rect 1868 1896 1876 1904
rect 1804 1876 1812 1884
rect 2092 1996 2100 2004
rect 2076 1976 2084 1984
rect 2140 1976 2148 1984
rect 2044 1956 2052 1964
rect 2060 1936 2068 1944
rect 2092 1956 2100 1964
rect 2012 1896 2020 1904
rect 2060 1896 2068 1904
rect 2108 1896 2116 1904
rect 2236 2016 2244 2024
rect 2220 1956 2228 1964
rect 2172 1936 2180 1944
rect 2220 1936 2228 1944
rect 2188 1896 2196 1904
rect 2364 2116 2372 2124
rect 2348 2076 2356 2084
rect 2380 2076 2388 2084
rect 2332 2016 2340 2024
rect 2412 2116 2420 2124
rect 2396 2036 2404 2044
rect 2556 2476 2564 2484
rect 2588 2476 2596 2484
rect 2524 2456 2532 2464
rect 2572 2456 2580 2464
rect 2572 2416 2580 2424
rect 2604 2456 2612 2464
rect 2572 2336 2580 2344
rect 2620 2436 2628 2444
rect 2700 2596 2708 2604
rect 2700 2576 2708 2584
rect 2748 2676 2756 2684
rect 2748 2576 2756 2584
rect 2700 2496 2708 2504
rect 2716 2456 2724 2464
rect 2700 2376 2708 2384
rect 2716 2376 2724 2384
rect 2508 2296 2516 2304
rect 2556 2296 2564 2304
rect 2636 2336 2644 2344
rect 2796 2836 2804 2844
rect 2860 2976 2868 2984
rect 2908 3036 2916 3044
rect 2956 3396 2964 3404
rect 2972 3376 2980 3384
rect 2972 3276 2980 3284
rect 2956 3256 2964 3264
rect 2956 3116 2964 3124
rect 2940 3056 2948 3064
rect 2924 2996 2932 3004
rect 2908 2976 2916 2984
rect 2924 2976 2932 2984
rect 2892 2956 2900 2964
rect 2876 2896 2884 2904
rect 2860 2776 2868 2784
rect 2860 2736 2868 2744
rect 2972 3076 2980 3084
rect 2972 2996 2980 3004
rect 2908 2896 2916 2904
rect 2924 2896 2932 2904
rect 2892 2856 2900 2864
rect 2892 2756 2900 2764
rect 2924 2816 2932 2824
rect 2796 2716 2804 2724
rect 2780 2696 2788 2704
rect 2828 2696 2836 2704
rect 2796 2676 2804 2684
rect 2844 2676 2852 2684
rect 2780 2656 2788 2664
rect 2828 2636 2836 2644
rect 2780 2556 2788 2564
rect 2796 2536 2804 2544
rect 2860 2636 2868 2644
rect 2844 2536 2852 2544
rect 2844 2516 2852 2524
rect 2876 2516 2884 2524
rect 2828 2476 2836 2484
rect 2860 2476 2868 2484
rect 2780 2456 2788 2464
rect 2620 2296 2628 2304
rect 2652 2296 2660 2304
rect 2684 2296 2692 2304
rect 2700 2296 2708 2304
rect 2508 2256 2516 2264
rect 2604 2256 2612 2264
rect 2668 2256 2676 2264
rect 2652 2236 2660 2244
rect 2492 2216 2500 2224
rect 2508 2196 2516 2204
rect 2476 2156 2484 2164
rect 2444 2116 2452 2124
rect 2572 2176 2580 2184
rect 2572 2136 2580 2144
rect 2428 2056 2436 2064
rect 2412 2016 2420 2024
rect 2444 2016 2452 2024
rect 2588 2116 2596 2124
rect 2556 2076 2564 2084
rect 2492 1976 2500 1984
rect 2332 1936 2340 1944
rect 2396 1936 2404 1944
rect 2508 1936 2516 1944
rect 2540 1936 2548 1944
rect 2236 1896 2244 1904
rect 2204 1876 2212 1884
rect 2268 1876 2276 1884
rect 2300 1876 2308 1884
rect 2044 1836 2052 1844
rect 2268 1836 2276 1844
rect 1772 1816 1780 1824
rect 1820 1816 1828 1824
rect 1724 1776 1732 1784
rect 1996 1776 2004 1784
rect 1708 1756 1716 1764
rect 1772 1756 1780 1764
rect 2012 1756 2020 1764
rect 1692 1736 1700 1744
rect 1644 1656 1652 1664
rect 1676 1696 1684 1704
rect 1708 1696 1716 1704
rect 1756 1696 1764 1704
rect 1692 1656 1700 1664
rect 1660 1576 1668 1584
rect 1692 1556 1700 1564
rect 1660 1516 1668 1524
rect 1788 1676 1796 1684
rect 1836 1656 1844 1664
rect 1884 1716 1892 1724
rect 1868 1696 1876 1704
rect 1932 1696 1940 1704
rect 1852 1636 1860 1644
rect 1820 1596 1828 1604
rect 1788 1496 1796 1504
rect 1724 1476 1732 1484
rect 1708 1456 1716 1464
rect 1660 1436 1668 1444
rect 1628 1376 1636 1384
rect 1676 1376 1684 1384
rect 1596 1336 1604 1344
rect 1324 1316 1332 1324
rect 1532 1316 1540 1324
rect 1564 1316 1572 1324
rect 1500 1296 1508 1304
rect 1532 1296 1540 1304
rect 1324 1276 1332 1284
rect 1548 1276 1556 1284
rect 1388 1256 1396 1264
rect 1340 1236 1348 1244
rect 1324 1196 1332 1204
rect 1276 1096 1284 1104
rect 1308 1096 1316 1104
rect 1244 1056 1252 1064
rect 1260 1036 1268 1044
rect 1228 896 1236 904
rect 1260 896 1268 904
rect 1308 996 1316 1004
rect 1660 1316 1668 1324
rect 1740 1376 1748 1384
rect 1692 1356 1700 1364
rect 1708 1356 1716 1364
rect 1852 1556 1860 1564
rect 1836 1516 1844 1524
rect 1916 1556 1924 1564
rect 1932 1536 1940 1544
rect 1836 1496 1844 1504
rect 1900 1496 1908 1504
rect 1916 1496 1924 1504
rect 1900 1456 1908 1464
rect 2060 1776 2068 1784
rect 2156 1776 2164 1784
rect 2124 1756 2132 1764
rect 2124 1736 2132 1744
rect 2156 1736 2164 1744
rect 2108 1716 2116 1724
rect 2236 1756 2244 1764
rect 2172 1716 2180 1724
rect 2220 1716 2228 1724
rect 2108 1696 2116 1704
rect 2156 1696 2164 1704
rect 2188 1696 2196 1704
rect 2044 1616 2052 1624
rect 2028 1576 2036 1584
rect 1996 1536 2004 1544
rect 1964 1476 1972 1484
rect 1980 1456 1988 1464
rect 2012 1456 2020 1464
rect 1692 1316 1700 1324
rect 1612 1296 1620 1304
rect 1676 1296 1684 1304
rect 1740 1296 1748 1304
rect 1788 1316 1796 1324
rect 1804 1296 1812 1304
rect 1964 1376 1972 1384
rect 1996 1376 2004 1384
rect 2012 1356 2020 1364
rect 1884 1316 1892 1324
rect 1644 1276 1652 1284
rect 1772 1276 1780 1284
rect 1612 1256 1620 1264
rect 1628 1256 1636 1264
rect 1836 1256 1844 1264
rect 1868 1256 1876 1264
rect 1596 1236 1604 1244
rect 1388 1216 1396 1224
rect 1404 1156 1412 1164
rect 1356 1116 1364 1124
rect 1452 1176 1460 1184
rect 1436 1156 1444 1164
rect 1566 1206 1574 1214
rect 1580 1206 1588 1214
rect 1594 1206 1602 1214
rect 1564 1176 1572 1184
rect 1516 1156 1524 1164
rect 1468 1136 1476 1144
rect 1500 1136 1508 1144
rect 1596 1136 1604 1144
rect 1468 1116 1476 1124
rect 1420 1096 1428 1104
rect 1452 1096 1460 1104
rect 1516 1096 1524 1104
rect 1612 1096 1620 1104
rect 1372 1076 1380 1084
rect 1740 1196 1748 1204
rect 1644 1176 1652 1184
rect 1756 1176 1764 1184
rect 1820 1176 1828 1184
rect 1820 1156 1828 1164
rect 1836 1156 1844 1164
rect 1724 1116 1732 1124
rect 1676 1096 1684 1104
rect 1660 1076 1668 1084
rect 1740 1096 1748 1104
rect 1724 1076 1732 1084
rect 1708 1056 1716 1064
rect 1724 1056 1732 1064
rect 1308 956 1316 964
rect 1228 776 1236 784
rect 1260 716 1268 724
rect 1228 696 1236 704
rect 1516 1016 1524 1024
rect 1404 976 1412 984
rect 1500 976 1508 984
rect 1708 976 1716 984
rect 1356 936 1364 944
rect 1388 916 1396 924
rect 1420 916 1428 924
rect 1340 896 1348 904
rect 1340 876 1348 884
rect 1372 876 1380 884
rect 1388 876 1396 884
rect 1324 836 1332 844
rect 1548 896 1556 904
rect 1452 856 1460 864
rect 1484 856 1492 864
rect 1660 896 1668 904
rect 1628 876 1636 884
rect 1612 856 1620 864
rect 1660 856 1668 864
rect 1692 856 1700 864
rect 1516 836 1524 844
rect 1564 836 1572 844
rect 1420 776 1428 784
rect 1308 756 1316 764
rect 1292 736 1300 744
rect 1276 676 1284 684
rect 1212 656 1220 664
rect 1292 656 1300 664
rect 924 636 932 644
rect 1004 636 1012 644
rect 1212 636 1220 644
rect 892 556 900 564
rect 892 516 900 524
rect 764 376 772 384
rect 764 356 772 364
rect 780 356 788 364
rect 732 316 740 324
rect 764 316 772 324
rect 716 296 724 304
rect 636 136 644 144
rect 652 116 660 124
rect 284 96 292 104
rect 332 96 340 104
rect 364 96 372 104
rect 508 96 516 104
rect 604 96 612 104
rect 684 96 692 104
rect 844 496 852 504
rect 860 456 868 464
rect 1004 596 1012 604
rect 1068 596 1076 604
rect 972 556 980 564
rect 956 516 964 524
rect 908 436 916 444
rect 828 416 836 424
rect 812 336 820 344
rect 844 396 852 404
rect 924 396 932 404
rect 908 316 916 324
rect 748 276 756 284
rect 780 276 788 284
rect 860 276 868 284
rect 876 256 884 264
rect 796 236 804 244
rect 1116 576 1124 584
rect 1372 736 1380 744
rect 1324 716 1332 724
rect 1420 716 1428 724
rect 1340 676 1348 684
rect 1388 656 1396 664
rect 1308 616 1316 624
rect 1356 616 1364 624
rect 1324 576 1332 584
rect 1228 556 1236 564
rect 1340 556 1348 564
rect 1132 536 1140 544
rect 1116 516 1124 524
rect 1004 476 1012 484
rect 988 456 996 464
rect 1052 456 1060 464
rect 1068 456 1076 464
rect 1068 436 1076 444
rect 1036 396 1044 404
rect 1020 376 1028 384
rect 988 336 996 344
rect 1020 336 1028 344
rect 1228 536 1236 544
rect 1292 536 1300 544
rect 1308 536 1316 544
rect 1164 516 1172 524
rect 1164 496 1172 504
rect 1116 416 1124 424
rect 1132 396 1140 404
rect 1324 516 1332 524
rect 1276 416 1284 424
rect 1356 536 1364 544
rect 1420 556 1428 564
rect 1566 806 1574 814
rect 1580 806 1588 814
rect 1594 806 1602 814
rect 1692 836 1700 844
rect 1548 776 1556 784
rect 1468 736 1476 744
rect 1564 736 1572 744
rect 1452 696 1460 704
rect 1516 656 1524 664
rect 1548 696 1556 704
rect 1724 896 1732 904
rect 1740 876 1748 884
rect 1772 1096 1780 1104
rect 1804 1036 1812 1044
rect 1820 1016 1828 1024
rect 2060 1516 2068 1524
rect 2124 1676 2132 1684
rect 2156 1676 2164 1684
rect 2156 1656 2164 1664
rect 2108 1516 2116 1524
rect 2092 1496 2100 1504
rect 2188 1596 2196 1604
rect 2172 1516 2180 1524
rect 2092 1456 2100 1464
rect 2140 1456 2148 1464
rect 2076 1436 2084 1444
rect 1948 1316 1956 1324
rect 2124 1396 2132 1404
rect 2108 1376 2116 1384
rect 2284 1676 2292 1684
rect 2332 1856 2340 1864
rect 2316 1696 2324 1704
rect 2364 1816 2372 1824
rect 2380 1796 2388 1804
rect 2364 1736 2372 1744
rect 2380 1696 2388 1704
rect 2348 1676 2356 1684
rect 2460 1896 2468 1904
rect 2492 1816 2500 1824
rect 2444 1796 2452 1804
rect 2476 1796 2484 1804
rect 2556 1816 2564 1824
rect 2604 2056 2612 2064
rect 2636 2076 2644 2084
rect 2636 1936 2644 1944
rect 2716 2236 2724 2244
rect 2764 2296 2772 2304
rect 2908 2716 2916 2724
rect 2956 2936 2964 2944
rect 2956 2816 2964 2824
rect 3052 3356 3060 3364
rect 3020 3296 3028 3304
rect 3004 3276 3012 3284
rect 3036 3256 3044 3264
rect 3228 3616 3236 3624
rect 3196 3536 3204 3544
rect 3244 3536 3252 3544
rect 3212 3516 3220 3524
rect 3244 3516 3252 3524
rect 3116 3476 3124 3484
rect 3212 3476 3220 3484
rect 3084 3456 3092 3464
rect 3132 3436 3140 3444
rect 3276 3696 3284 3704
rect 3308 3676 3316 3684
rect 3356 3736 3364 3744
rect 3340 3696 3348 3704
rect 3516 4156 3524 4164
rect 3548 4156 3556 4164
rect 3548 4136 3556 4144
rect 3692 4336 3700 4344
rect 3660 4296 3668 4304
rect 3676 4296 3684 4304
rect 3612 4176 3620 4184
rect 3644 4216 3652 4224
rect 3628 4136 3636 4144
rect 3532 4016 3540 4024
rect 3404 3896 3412 3904
rect 3436 3896 3444 3904
rect 3484 3896 3492 3904
rect 3436 3836 3444 3844
rect 3420 3816 3428 3824
rect 3452 3816 3460 3824
rect 3436 3756 3444 3764
rect 3516 3896 3524 3904
rect 3580 3976 3588 3984
rect 3548 3916 3556 3924
rect 3596 3936 3604 3944
rect 3564 3876 3572 3884
rect 3580 3856 3588 3864
rect 3596 3836 3604 3844
rect 3548 3776 3556 3784
rect 3804 4496 3812 4504
rect 3740 4456 3748 4464
rect 3868 4396 3876 4404
rect 3820 4336 3828 4344
rect 3724 4296 3732 4304
rect 3740 4296 3748 4304
rect 3772 4296 3780 4304
rect 3724 4276 3732 4284
rect 3724 4256 3732 4264
rect 3708 4236 3716 4244
rect 3788 4276 3796 4284
rect 3804 4276 3812 4284
rect 3820 4256 3828 4264
rect 3884 4276 3892 4284
rect 3948 4496 3956 4504
rect 3916 4436 3924 4444
rect 3948 4476 3956 4484
rect 3932 4396 3940 4404
rect 3996 4436 4004 4444
rect 3996 4336 4004 4344
rect 4460 4936 4468 4944
rect 4444 4896 4452 4904
rect 4412 4876 4420 4884
rect 4316 4776 4324 4784
rect 4252 4756 4260 4764
rect 4300 4756 4308 4764
rect 4364 4756 4372 4764
rect 4380 4756 4388 4764
rect 4316 4736 4324 4744
rect 4380 4736 4388 4744
rect 4396 4736 4404 4744
rect 4204 4716 4212 4724
rect 4204 4676 4212 4684
rect 4236 4676 4244 4684
rect 4412 4716 4420 4724
rect 4332 4696 4340 4704
rect 4380 4676 4388 4684
rect 4412 4676 4420 4684
rect 4268 4656 4276 4664
rect 4252 4636 4260 4644
rect 4284 4596 4292 4604
rect 4412 4656 4420 4664
rect 4428 4656 4436 4664
rect 4396 4636 4404 4644
rect 4236 4576 4244 4584
rect 4092 4556 4100 4564
rect 4156 4556 4164 4564
rect 4300 4556 4308 4564
rect 4092 4536 4100 4544
rect 4124 4536 4132 4544
rect 4188 4536 4196 4544
rect 4252 4536 4260 4544
rect 4284 4536 4292 4544
rect 4140 4496 4148 4504
rect 4124 4456 4132 4464
rect 4076 4436 4084 4444
rect 4044 4336 4052 4344
rect 4108 4336 4116 4344
rect 3852 4236 3860 4244
rect 3900 4236 3908 4244
rect 3772 4156 3780 4164
rect 3740 4136 3748 4144
rect 3628 4116 3636 4124
rect 3676 3976 3684 3984
rect 3692 3976 3700 3984
rect 3660 3936 3668 3944
rect 3628 3896 3636 3904
rect 3740 4076 3748 4084
rect 3820 4136 3828 4144
rect 3788 4116 3796 4124
rect 3756 4036 3764 4044
rect 3932 4296 3940 4304
rect 3932 4276 3940 4284
rect 3804 4076 3812 4084
rect 3804 4056 3812 4064
rect 3740 3956 3748 3964
rect 3788 3956 3796 3964
rect 3724 3916 3732 3924
rect 3772 3916 3780 3924
rect 3612 3816 3620 3824
rect 3708 3836 3716 3844
rect 3692 3816 3700 3824
rect 3756 3816 3764 3824
rect 3628 3756 3636 3764
rect 3404 3636 3412 3644
rect 3356 3596 3364 3604
rect 3324 3576 3332 3584
rect 3308 3536 3316 3544
rect 3404 3536 3412 3544
rect 3292 3516 3300 3524
rect 3260 3496 3268 3504
rect 3292 3496 3300 3504
rect 3276 3436 3284 3444
rect 3212 3416 3220 3424
rect 3244 3416 3252 3424
rect 3260 3416 3268 3424
rect 3118 3406 3126 3414
rect 3132 3406 3140 3414
rect 3146 3406 3154 3414
rect 3196 3376 3204 3384
rect 3228 3356 3236 3364
rect 3148 3336 3156 3344
rect 3180 3316 3188 3324
rect 3228 3316 3236 3324
rect 3164 3296 3172 3304
rect 3356 3516 3364 3524
rect 3324 3496 3332 3504
rect 3340 3456 3348 3464
rect 3324 3416 3332 3424
rect 3340 3416 3348 3424
rect 3260 3336 3268 3344
rect 3260 3316 3268 3324
rect 3132 3256 3140 3264
rect 3212 3276 3220 3284
rect 3308 3316 3316 3324
rect 3292 3256 3300 3264
rect 3388 3476 3396 3484
rect 3356 3356 3364 3364
rect 3372 3356 3380 3364
rect 3356 3336 3364 3344
rect 3324 3296 3332 3304
rect 3068 3156 3076 3164
rect 3196 3156 3204 3164
rect 3260 3156 3268 3164
rect 3036 3116 3044 3124
rect 3004 3096 3012 3104
rect 3020 3076 3028 3084
rect 3004 3016 3012 3024
rect 2988 2956 2996 2964
rect 3004 2956 3012 2964
rect 3004 2936 3012 2944
rect 2988 2916 2996 2924
rect 2988 2896 2996 2904
rect 3004 2896 3012 2904
rect 3036 2996 3044 3004
rect 3036 2976 3044 2984
rect 3180 3136 3188 3144
rect 3132 3116 3140 3124
rect 3084 3096 3092 3104
rect 3164 3076 3172 3084
rect 3164 3036 3172 3044
rect 3118 3006 3126 3014
rect 3132 3006 3140 3014
rect 3146 3006 3154 3014
rect 3228 3136 3236 3144
rect 3212 3056 3220 3064
rect 3180 2996 3188 3004
rect 3100 2976 3108 2984
rect 3212 2976 3220 2984
rect 3196 2956 3204 2964
rect 3068 2936 3076 2944
rect 3148 2936 3156 2944
rect 3196 2936 3204 2944
rect 3212 2936 3220 2944
rect 3052 2916 3060 2924
rect 3036 2896 3044 2904
rect 3020 2876 3028 2884
rect 3004 2836 3012 2844
rect 2988 2816 2996 2824
rect 3020 2716 3028 2724
rect 3020 2676 3028 2684
rect 2940 2636 2948 2644
rect 2988 2636 2996 2644
rect 2972 2616 2980 2624
rect 2940 2596 2948 2604
rect 2924 2516 2932 2524
rect 3084 2896 3092 2904
rect 3180 2896 3188 2904
rect 3212 2896 3220 2904
rect 3068 2876 3076 2884
rect 3052 2856 3060 2864
rect 3068 2856 3076 2864
rect 3052 2656 3060 2664
rect 3084 2836 3092 2844
rect 3100 2836 3108 2844
rect 3084 2816 3092 2824
rect 3116 2816 3124 2824
rect 3084 2716 3092 2724
rect 3100 2716 3108 2724
rect 3068 2636 3076 2644
rect 2988 2556 2996 2564
rect 2988 2516 2996 2524
rect 2908 2496 2916 2504
rect 3020 2496 3028 2504
rect 2940 2476 2948 2484
rect 3020 2476 3028 2484
rect 2924 2436 2932 2444
rect 2844 2396 2852 2404
rect 2892 2396 2900 2404
rect 2924 2396 2932 2404
rect 2796 2316 2804 2324
rect 2812 2316 2820 2324
rect 2892 2316 2900 2324
rect 2860 2296 2868 2304
rect 2876 2296 2884 2304
rect 2844 2276 2852 2284
rect 2780 2256 2788 2264
rect 2828 2256 2836 2264
rect 2812 2236 2820 2244
rect 2812 2136 2820 2144
rect 2780 2116 2788 2124
rect 2732 2076 2740 2084
rect 2796 2056 2804 2064
rect 2700 2036 2708 2044
rect 2684 2016 2692 2024
rect 2588 1856 2596 1864
rect 2716 2016 2724 2024
rect 2764 1956 2772 1964
rect 2812 1956 2820 1964
rect 2732 1936 2740 1944
rect 2796 1936 2804 1944
rect 2684 1896 2692 1904
rect 2700 1876 2708 1884
rect 2620 1816 2628 1824
rect 2572 1796 2580 1804
rect 2636 1796 2644 1804
rect 2476 1776 2484 1784
rect 2444 1716 2452 1724
rect 2476 1716 2484 1724
rect 2412 1676 2420 1684
rect 2428 1676 2436 1684
rect 2588 1736 2596 1744
rect 2604 1716 2612 1724
rect 2460 1696 2468 1704
rect 2524 1696 2532 1704
rect 2540 1676 2548 1684
rect 2572 1676 2580 1684
rect 2748 1896 2756 1904
rect 2764 1896 2772 1904
rect 2732 1836 2740 1844
rect 2716 1756 2724 1764
rect 2732 1756 2740 1764
rect 2700 1736 2708 1744
rect 2668 1716 2676 1724
rect 2620 1656 2628 1664
rect 2636 1656 2644 1664
rect 2380 1636 2388 1644
rect 2396 1636 2404 1644
rect 2476 1636 2484 1644
rect 2380 1596 2388 1604
rect 2748 1736 2756 1744
rect 2716 1696 2724 1704
rect 2748 1696 2756 1704
rect 2668 1616 2676 1624
rect 2220 1576 2228 1584
rect 2268 1576 2276 1584
rect 2332 1576 2340 1584
rect 2460 1576 2468 1584
rect 2204 1496 2212 1504
rect 2188 1456 2196 1464
rect 2204 1436 2212 1444
rect 2396 1556 2404 1564
rect 2284 1536 2292 1544
rect 2236 1436 2244 1444
rect 2252 1396 2260 1404
rect 2268 1376 2276 1384
rect 2172 1356 2180 1364
rect 2092 1336 2100 1344
rect 2188 1336 2196 1344
rect 2060 1316 2068 1324
rect 2140 1316 2148 1324
rect 1932 1196 1940 1204
rect 1964 1276 1972 1284
rect 1948 1176 1956 1184
rect 1900 1136 1908 1144
rect 1948 1136 1956 1144
rect 1868 1096 1876 1104
rect 1884 1096 1892 1104
rect 1852 1016 1860 1024
rect 1964 1076 1972 1084
rect 1900 1056 1908 1064
rect 1772 956 1780 964
rect 1820 956 1828 964
rect 1836 956 1844 964
rect 1788 896 1796 904
rect 1836 936 1844 944
rect 1884 916 1892 924
rect 1836 896 1844 904
rect 1804 876 1812 884
rect 1756 756 1764 764
rect 1804 796 1812 804
rect 1772 696 1780 704
rect 1740 676 1748 684
rect 1596 616 1604 624
rect 1612 576 1620 584
rect 1676 576 1684 584
rect 1532 556 1540 564
rect 1340 456 1348 464
rect 1372 456 1380 464
rect 1436 536 1444 544
rect 1420 456 1428 464
rect 1388 436 1396 444
rect 1404 436 1412 444
rect 1244 376 1252 384
rect 1084 356 1092 364
rect 1196 356 1204 364
rect 1372 356 1380 364
rect 1068 336 1076 344
rect 1084 336 1092 344
rect 1116 336 1124 344
rect 1180 336 1188 344
rect 1260 336 1268 344
rect 1308 336 1316 344
rect 1324 336 1332 344
rect 1388 336 1396 344
rect 988 316 996 324
rect 1004 316 1012 324
rect 1212 316 1220 324
rect 956 296 964 304
rect 972 296 980 304
rect 924 236 932 244
rect 1132 296 1140 304
rect 1100 276 1108 284
rect 1052 256 1060 264
rect 908 216 916 224
rect 972 216 980 224
rect 860 196 868 204
rect 1020 236 1028 244
rect 1004 216 1012 224
rect 796 156 804 164
rect 812 156 820 164
rect 988 156 996 164
rect 1004 156 1012 164
rect 732 136 740 144
rect 748 116 756 124
rect 780 116 788 124
rect 860 116 868 124
rect 940 116 948 124
rect 732 96 740 104
rect 764 96 772 104
rect 620 76 628 84
rect 1116 256 1124 264
rect 1196 296 1204 304
rect 1244 296 1252 304
rect 1244 276 1252 284
rect 1340 316 1348 324
rect 1484 516 1492 524
rect 1500 516 1508 524
rect 1468 436 1476 444
rect 1500 396 1508 404
rect 1548 516 1556 524
rect 1612 516 1620 524
rect 1868 836 1876 844
rect 1948 1036 1956 1044
rect 2044 1296 2052 1304
rect 2140 1296 2148 1304
rect 2156 1296 2164 1304
rect 2012 1256 2020 1264
rect 2028 1256 2036 1264
rect 1996 1136 2004 1144
rect 2076 1216 2084 1224
rect 2140 1216 2148 1224
rect 2076 1136 2084 1144
rect 2124 1136 2132 1144
rect 2140 1136 2148 1144
rect 1996 1116 2004 1124
rect 2012 1116 2020 1124
rect 2012 1076 2020 1084
rect 1980 976 1988 984
rect 1964 956 1972 964
rect 1948 916 1956 924
rect 1948 896 1956 904
rect 1932 876 1940 884
rect 1884 776 1892 784
rect 1868 756 1876 764
rect 1820 736 1828 744
rect 1820 716 1828 724
rect 1852 716 1860 724
rect 1836 676 1844 684
rect 1884 736 1892 744
rect 1900 676 1908 684
rect 1916 596 1924 604
rect 1948 836 1956 844
rect 1964 836 1972 844
rect 1996 896 2004 904
rect 2252 1316 2260 1324
rect 2236 1296 2244 1304
rect 2236 1276 2244 1284
rect 2204 1236 2212 1244
rect 2188 1196 2196 1204
rect 2172 1176 2180 1184
rect 2092 1116 2100 1124
rect 2140 1116 2148 1124
rect 2156 1116 2164 1124
rect 2140 1076 2148 1084
rect 2060 996 2068 1004
rect 2028 956 2036 964
rect 2028 916 2036 924
rect 2044 856 2052 864
rect 2076 956 2084 964
rect 2092 936 2100 944
rect 2108 856 2116 864
rect 2012 796 2020 804
rect 2028 796 2036 804
rect 1948 636 1956 644
rect 1980 696 1988 704
rect 1964 576 1972 584
rect 1772 536 1780 544
rect 1676 516 1684 524
rect 1692 496 1700 504
rect 1740 496 1748 504
rect 1660 476 1668 484
rect 1724 476 1732 484
rect 1788 496 1796 504
rect 1772 476 1780 484
rect 1836 516 1844 524
rect 1628 456 1636 464
rect 1708 456 1716 464
rect 1756 456 1764 464
rect 1820 456 1828 464
rect 1566 406 1574 414
rect 1580 406 1588 414
rect 1594 406 1602 414
rect 1644 396 1652 404
rect 1692 376 1700 384
rect 1484 356 1492 364
rect 1612 356 1620 364
rect 1676 356 1684 364
rect 1516 336 1524 344
rect 1324 296 1332 304
rect 1372 296 1380 304
rect 1276 276 1284 284
rect 1308 276 1316 284
rect 1324 276 1332 284
rect 1260 236 1268 244
rect 1276 236 1284 244
rect 1148 216 1156 224
rect 1228 216 1236 224
rect 1260 216 1268 224
rect 1164 176 1172 184
rect 1148 156 1156 164
rect 1388 236 1396 244
rect 1436 296 1444 304
rect 1484 296 1492 304
rect 1452 256 1460 264
rect 1500 216 1508 224
rect 1420 196 1428 204
rect 1484 196 1492 204
rect 1292 156 1300 164
rect 1372 156 1380 164
rect 1436 156 1444 164
rect 1500 156 1508 164
rect 1228 136 1236 144
rect 1308 136 1316 144
rect 1340 136 1348 144
rect 1404 136 1412 144
rect 1436 136 1444 144
rect 1244 116 1252 124
rect 1100 96 1108 104
rect 876 76 884 84
rect 908 76 916 84
rect 956 76 964 84
rect 1068 76 1076 84
rect 1116 76 1124 84
rect 284 56 292 64
rect 844 56 852 64
rect 924 56 932 64
rect 1356 96 1364 104
rect 1388 96 1396 104
rect 1564 296 1572 304
rect 1628 336 1636 344
rect 1804 416 1812 424
rect 1740 316 1748 324
rect 1788 296 1796 304
rect 1724 276 1732 284
rect 1692 256 1700 264
rect 1724 256 1732 264
rect 1724 236 1732 244
rect 1596 216 1604 224
rect 1564 196 1572 204
rect 1788 216 1796 224
rect 1740 196 1748 204
rect 1916 516 1924 524
rect 1996 616 2004 624
rect 2028 636 2036 644
rect 2012 576 2020 584
rect 2108 836 2116 844
rect 2092 736 2100 744
rect 2060 716 2068 724
rect 2108 676 2116 684
rect 2220 1196 2228 1204
rect 2268 1236 2276 1244
rect 2332 1516 2340 1524
rect 2716 1616 2724 1624
rect 2732 1556 2740 1564
rect 2444 1536 2452 1544
rect 2700 1536 2708 1544
rect 2716 1536 2724 1544
rect 2380 1516 2388 1524
rect 2428 1516 2436 1524
rect 2300 1496 2308 1504
rect 2364 1496 2372 1504
rect 2316 1476 2324 1484
rect 2540 1496 2548 1504
rect 2588 1496 2596 1504
rect 2412 1476 2420 1484
rect 2316 1376 2324 1384
rect 2332 1376 2340 1384
rect 2364 1376 2372 1384
rect 2300 1316 2308 1324
rect 2316 1276 2324 1284
rect 2300 1236 2308 1244
rect 2252 1136 2260 1144
rect 2220 1116 2228 1124
rect 2252 1116 2260 1124
rect 2172 1076 2180 1084
rect 2172 1036 2180 1044
rect 2348 1316 2356 1324
rect 2412 1436 2420 1444
rect 2396 1336 2404 1344
rect 2396 1316 2404 1324
rect 2652 1496 2660 1504
rect 2700 1496 2708 1504
rect 2812 1816 2820 1824
rect 2812 1776 2820 1784
rect 2796 1756 2804 1764
rect 2812 1736 2820 1744
rect 2796 1696 2804 1704
rect 2780 1536 2788 1544
rect 2764 1496 2772 1504
rect 2492 1476 2500 1484
rect 2556 1476 2564 1484
rect 2588 1476 2596 1484
rect 2620 1476 2628 1484
rect 2652 1476 2660 1484
rect 2748 1476 2756 1484
rect 2476 1436 2484 1444
rect 2508 1436 2516 1444
rect 2492 1416 2500 1424
rect 2476 1396 2484 1404
rect 2556 1416 2564 1424
rect 2540 1396 2548 1404
rect 2524 1356 2532 1364
rect 2508 1336 2516 1344
rect 2444 1316 2452 1324
rect 2476 1316 2484 1324
rect 2412 1276 2420 1284
rect 2396 1216 2404 1224
rect 2428 1196 2436 1204
rect 2348 1176 2356 1184
rect 2396 1156 2404 1164
rect 2348 1136 2356 1144
rect 2332 1116 2340 1124
rect 2300 1076 2308 1084
rect 2348 1056 2356 1064
rect 2380 1076 2388 1084
rect 2268 1016 2276 1024
rect 2236 996 2244 1004
rect 2332 976 2340 984
rect 2284 936 2292 944
rect 2220 916 2228 924
rect 2268 916 2276 924
rect 2300 916 2308 924
rect 2204 896 2212 904
rect 2188 876 2196 884
rect 2332 876 2340 884
rect 2188 856 2196 864
rect 2172 836 2180 844
rect 2188 816 2196 824
rect 2156 776 2164 784
rect 2204 756 2212 764
rect 2140 736 2148 744
rect 2188 696 2196 704
rect 2172 676 2180 684
rect 2156 656 2164 664
rect 2140 616 2148 624
rect 2076 556 2084 564
rect 2092 556 2100 564
rect 1884 476 1892 484
rect 1932 476 1940 484
rect 1980 476 1988 484
rect 2028 476 2036 484
rect 1932 456 1940 464
rect 1852 436 1860 444
rect 1900 436 1908 444
rect 1836 396 1844 404
rect 2172 536 2180 544
rect 2380 1036 2388 1044
rect 2556 1336 2564 1344
rect 2588 1296 2596 1304
rect 2524 1256 2532 1264
rect 2572 1256 2580 1264
rect 2508 1216 2516 1224
rect 2492 1196 2500 1204
rect 2444 1136 2452 1144
rect 2428 1116 2436 1124
rect 2428 1076 2436 1084
rect 2412 976 2420 984
rect 2444 1036 2452 1044
rect 2460 916 2468 924
rect 2476 916 2484 924
rect 2396 896 2404 904
rect 2620 1296 2628 1304
rect 2620 1256 2628 1264
rect 2604 1176 2612 1184
rect 2684 1436 2692 1444
rect 2716 1456 2724 1464
rect 2700 1376 2708 1384
rect 2668 1356 2676 1364
rect 2716 1316 2724 1324
rect 2700 1216 2708 1224
rect 2620 1156 2628 1164
rect 2636 1156 2644 1164
rect 2572 1136 2580 1144
rect 2588 1116 2596 1124
rect 2508 1096 2516 1104
rect 2572 1076 2580 1084
rect 2540 1056 2548 1064
rect 2524 1016 2532 1024
rect 2556 996 2564 1004
rect 2540 976 2548 984
rect 2524 896 2532 904
rect 2396 876 2404 884
rect 2492 876 2500 884
rect 2364 816 2372 824
rect 2380 776 2388 784
rect 2460 776 2468 784
rect 2348 756 2356 764
rect 2428 756 2436 764
rect 2252 736 2260 744
rect 2444 736 2452 744
rect 2236 716 2244 724
rect 2364 716 2372 724
rect 2412 716 2420 724
rect 2220 696 2228 704
rect 2284 696 2292 704
rect 2252 576 2260 584
rect 2492 736 2500 744
rect 2540 876 2548 884
rect 2700 1176 2708 1184
rect 2668 1156 2676 1164
rect 2652 1116 2660 1124
rect 2764 1456 2772 1464
rect 2764 1316 2772 1324
rect 2812 1676 2820 1684
rect 2844 2076 2852 2084
rect 2844 2056 2852 2064
rect 2844 1936 2852 1944
rect 2908 2276 2916 2284
rect 2876 2236 2884 2244
rect 2972 2416 2980 2424
rect 3004 2416 3012 2424
rect 2956 2316 2964 2324
rect 2972 2316 2980 2324
rect 3004 2316 3012 2324
rect 2940 2296 2948 2304
rect 2924 2196 2932 2204
rect 2876 2176 2884 2184
rect 2892 2156 2900 2164
rect 2956 2276 2964 2284
rect 3196 2816 3204 2824
rect 3212 2816 3220 2824
rect 3180 2776 3188 2784
rect 3212 2776 3220 2784
rect 3164 2756 3172 2764
rect 3180 2756 3188 2764
rect 3196 2736 3204 2744
rect 3244 3096 3252 3104
rect 3276 3056 3284 3064
rect 3260 2996 3268 3004
rect 3276 2996 3284 3004
rect 3244 2956 3252 2964
rect 3308 3096 3316 3104
rect 3436 3636 3444 3644
rect 3500 3736 3508 3744
rect 3468 3696 3476 3704
rect 3484 3696 3492 3704
rect 3468 3556 3476 3564
rect 3452 3516 3460 3524
rect 3500 3676 3508 3684
rect 3500 3636 3508 3644
rect 3484 3536 3492 3544
rect 3484 3476 3492 3484
rect 3452 3376 3460 3384
rect 3420 3356 3428 3364
rect 3452 3356 3460 3364
rect 3420 3316 3428 3324
rect 3372 3296 3380 3304
rect 3388 3276 3396 3284
rect 3420 3276 3428 3284
rect 3420 3256 3428 3264
rect 3404 3236 3412 3244
rect 3388 3216 3396 3224
rect 3372 3176 3380 3184
rect 3372 3156 3380 3164
rect 3356 3036 3364 3044
rect 3324 2976 3332 2984
rect 3308 2956 3316 2964
rect 3308 2936 3316 2944
rect 3292 2916 3300 2924
rect 3292 2896 3300 2904
rect 3276 2856 3284 2864
rect 3228 2756 3236 2764
rect 3164 2716 3172 2724
rect 3212 2716 3220 2724
rect 3212 2696 3220 2704
rect 3180 2636 3188 2644
rect 3196 2636 3204 2644
rect 3118 2606 3126 2614
rect 3132 2606 3140 2614
rect 3146 2606 3154 2614
rect 3244 2696 3252 2704
rect 3228 2616 3236 2624
rect 3148 2576 3156 2584
rect 3180 2576 3188 2584
rect 3164 2556 3172 2564
rect 3164 2516 3172 2524
rect 3196 2516 3204 2524
rect 3068 2436 3076 2444
rect 3084 2436 3092 2444
rect 3100 2416 3108 2424
rect 3084 2316 3092 2324
rect 3020 2296 3028 2304
rect 3036 2296 3044 2304
rect 2988 2276 2996 2284
rect 2972 2236 2980 2244
rect 2988 2236 2996 2244
rect 3020 2276 3028 2284
rect 2956 2156 2964 2164
rect 2940 2136 2948 2144
rect 2908 2076 2916 2084
rect 2892 2036 2900 2044
rect 3052 2276 3060 2284
rect 3116 2376 3124 2384
rect 3276 2676 3284 2684
rect 3324 2916 3332 2924
rect 3356 2916 3364 2924
rect 3356 2776 3364 2784
rect 3356 2736 3364 2744
rect 3356 2696 3364 2704
rect 3308 2676 3316 2684
rect 3436 3196 3444 3204
rect 3484 3316 3492 3324
rect 3532 3736 3540 3744
rect 3612 3736 3620 3744
rect 3708 3736 3716 3744
rect 3532 3696 3540 3704
rect 3548 3696 3556 3704
rect 3532 3616 3540 3624
rect 3516 3476 3524 3484
rect 3516 3456 3524 3464
rect 3516 3376 3524 3384
rect 3516 3316 3524 3324
rect 3500 3176 3508 3184
rect 3468 3156 3476 3164
rect 3468 3136 3476 3144
rect 3420 3116 3428 3124
rect 3388 3016 3396 3024
rect 3436 3096 3444 3104
rect 3676 3696 3684 3704
rect 3580 3676 3588 3684
rect 3628 3576 3636 3584
rect 3596 3536 3604 3544
rect 3564 3516 3572 3524
rect 3548 3496 3556 3504
rect 3548 3456 3556 3464
rect 3692 3536 3700 3544
rect 3628 3476 3636 3484
rect 3612 3436 3620 3444
rect 3564 3316 3572 3324
rect 3532 3256 3540 3264
rect 3548 3176 3556 3184
rect 3580 3296 3588 3304
rect 3660 3476 3668 3484
rect 3676 3456 3684 3464
rect 3644 3416 3652 3424
rect 3676 3416 3684 3424
rect 3660 3376 3668 3384
rect 3628 3296 3636 3304
rect 3596 3276 3604 3284
rect 3612 3276 3620 3284
rect 3580 3256 3588 3264
rect 3532 3136 3540 3144
rect 3500 3076 3508 3084
rect 3420 3056 3428 3064
rect 3452 3056 3460 3064
rect 3468 3036 3476 3044
rect 3436 3016 3444 3024
rect 3452 3016 3460 3024
rect 3404 2996 3412 3004
rect 3420 2996 3428 3004
rect 3404 2976 3412 2984
rect 3452 2916 3460 2924
rect 3484 2936 3492 2944
rect 3484 2916 3492 2924
rect 3452 2896 3460 2904
rect 3468 2896 3476 2904
rect 3420 2876 3428 2884
rect 3404 2836 3412 2844
rect 3388 2796 3396 2804
rect 3388 2676 3396 2684
rect 3324 2636 3332 2644
rect 3340 2636 3348 2644
rect 3372 2636 3380 2644
rect 3276 2616 3284 2624
rect 3292 2616 3300 2624
rect 3260 2596 3268 2604
rect 3260 2576 3268 2584
rect 3260 2536 3268 2544
rect 3244 2496 3252 2504
rect 3212 2476 3220 2484
rect 3228 2476 3236 2484
rect 3148 2376 3156 2384
rect 3132 2356 3140 2364
rect 3260 2416 3268 2424
rect 3356 2616 3364 2624
rect 3404 2616 3412 2624
rect 3356 2556 3364 2564
rect 3324 2496 3332 2504
rect 3340 2476 3348 2484
rect 3308 2456 3316 2464
rect 3292 2416 3300 2424
rect 3276 2356 3284 2364
rect 3340 2356 3348 2364
rect 3180 2316 3188 2324
rect 3212 2316 3220 2324
rect 3260 2316 3268 2324
rect 3292 2316 3300 2324
rect 3324 2316 3332 2324
rect 3148 2296 3156 2304
rect 3068 2256 3076 2264
rect 3100 2256 3108 2264
rect 3196 2296 3204 2304
rect 3164 2256 3172 2264
rect 3196 2256 3204 2264
rect 3084 2236 3092 2244
rect 3148 2236 3156 2244
rect 3036 2216 3044 2224
rect 3036 2196 3044 2204
rect 3068 2156 3076 2164
rect 3052 2136 3060 2144
rect 3036 2036 3044 2044
rect 3004 2016 3012 2024
rect 3020 2016 3028 2024
rect 3180 2216 3188 2224
rect 3118 2206 3126 2214
rect 3132 2206 3140 2214
rect 3146 2206 3154 2214
rect 3388 2536 3396 2544
rect 3468 2756 3476 2764
rect 3516 3056 3524 3064
rect 3532 3036 3540 3044
rect 3516 2976 3524 2984
rect 3596 3096 3604 3104
rect 3628 3136 3636 3144
rect 3644 3116 3652 3124
rect 3644 3076 3652 3084
rect 3564 3036 3572 3044
rect 3612 3016 3620 3024
rect 3596 2976 3604 2984
rect 3548 2956 3556 2964
rect 3564 2936 3572 2944
rect 3516 2896 3524 2904
rect 3500 2876 3508 2884
rect 3516 2816 3524 2824
rect 3548 2816 3556 2824
rect 3532 2796 3540 2804
rect 3612 2936 3620 2944
rect 3580 2836 3588 2844
rect 3596 2836 3604 2844
rect 3628 2796 3636 2804
rect 3580 2776 3588 2784
rect 3596 2776 3604 2784
rect 3564 2756 3572 2764
rect 3484 2736 3492 2744
rect 3548 2736 3556 2744
rect 3580 2736 3588 2744
rect 3484 2716 3492 2724
rect 3468 2676 3476 2684
rect 3452 2636 3460 2644
rect 3468 2636 3476 2644
rect 3436 2616 3444 2624
rect 3468 2576 3476 2584
rect 3532 2716 3540 2724
rect 3516 2676 3524 2684
rect 3420 2536 3428 2544
rect 3452 2536 3460 2544
rect 3244 2296 3252 2304
rect 3260 2296 3268 2304
rect 3308 2296 3316 2304
rect 3340 2296 3348 2304
rect 3356 2296 3364 2304
rect 3244 2256 3252 2264
rect 3276 2256 3284 2264
rect 3212 2196 3220 2204
rect 3228 2176 3236 2184
rect 3260 2216 3268 2224
rect 3276 2196 3284 2204
rect 3260 2176 3268 2184
rect 3228 2136 3236 2144
rect 3132 2076 3140 2084
rect 3148 2076 3156 2084
rect 3100 2036 3108 2044
rect 3132 2036 3140 2044
rect 3100 2016 3108 2024
rect 2940 1976 2948 1984
rect 3036 1976 3044 1984
rect 3052 1976 3060 1984
rect 3068 1976 3076 1984
rect 2924 1956 2932 1964
rect 2892 1916 2900 1924
rect 2876 1896 2884 1904
rect 2860 1876 2868 1884
rect 2924 1836 2932 1844
rect 2876 1796 2884 1804
rect 2892 1796 2900 1804
rect 2844 1776 2852 1784
rect 2812 1636 2820 1644
rect 2860 1676 2868 1684
rect 2844 1596 2852 1604
rect 2972 1956 2980 1964
rect 2956 1916 2964 1924
rect 2988 1916 2996 1924
rect 2972 1896 2980 1904
rect 3004 1896 3012 1904
rect 3052 1916 3060 1924
rect 3036 1896 3044 1904
rect 2988 1876 2996 1884
rect 2972 1856 2980 1864
rect 2956 1796 2964 1804
rect 2892 1776 2900 1784
rect 2940 1776 2948 1784
rect 2908 1756 2916 1764
rect 2876 1596 2884 1604
rect 2860 1576 2868 1584
rect 2828 1536 2836 1544
rect 2860 1536 2868 1544
rect 2892 1536 2900 1544
rect 2812 1516 2820 1524
rect 2828 1516 2836 1524
rect 2924 1676 2932 1684
rect 2972 1656 2980 1664
rect 2924 1616 2932 1624
rect 2940 1616 2948 1624
rect 2924 1556 2932 1564
rect 2796 1456 2804 1464
rect 2876 1456 2884 1464
rect 2812 1436 2820 1444
rect 2812 1396 2820 1404
rect 2844 1376 2852 1384
rect 2876 1416 2884 1424
rect 2860 1336 2868 1344
rect 2876 1316 2884 1324
rect 2780 1296 2788 1304
rect 2812 1296 2820 1304
rect 2748 1256 2756 1264
rect 2796 1236 2804 1244
rect 3068 1896 3076 1904
rect 3036 1856 3044 1864
rect 3020 1796 3028 1804
rect 3004 1776 3012 1784
rect 3020 1696 3028 1704
rect 3164 1976 3172 1984
rect 3196 2076 3204 2084
rect 3244 2076 3252 2084
rect 3196 2056 3204 2064
rect 3228 2056 3236 2064
rect 3180 1956 3188 1964
rect 3196 1956 3204 1964
rect 3212 1956 3220 1964
rect 3100 1916 3108 1924
rect 3100 1896 3108 1904
rect 3180 1896 3188 1904
rect 3084 1836 3092 1844
rect 3116 1836 3124 1844
rect 3068 1816 3076 1824
rect 3052 1736 3060 1744
rect 3118 1806 3126 1814
rect 3132 1806 3140 1814
rect 3146 1806 3154 1814
rect 3116 1776 3124 1784
rect 3100 1756 3108 1764
rect 3036 1676 3044 1684
rect 3020 1636 3028 1644
rect 3100 1676 3108 1684
rect 2988 1576 2996 1584
rect 3068 1576 3076 1584
rect 2956 1556 2964 1564
rect 3020 1556 3028 1564
rect 3068 1556 3076 1564
rect 3212 1916 3220 1924
rect 3308 2216 3316 2224
rect 3356 2276 3364 2284
rect 3404 2496 3412 2504
rect 3484 2536 3492 2544
rect 3452 2456 3460 2464
rect 3468 2456 3476 2464
rect 3500 2476 3508 2484
rect 3468 2396 3476 2404
rect 3484 2396 3492 2404
rect 3404 2376 3412 2384
rect 3388 2316 3396 2324
rect 3372 2176 3380 2184
rect 3308 2136 3316 2144
rect 3340 2136 3348 2144
rect 3372 2136 3380 2144
rect 3356 2096 3364 2104
rect 3292 2076 3300 2084
rect 3340 2076 3348 2084
rect 3276 2056 3284 2064
rect 3260 1976 3268 1984
rect 3276 1976 3284 1984
rect 3292 1916 3300 1924
rect 3276 1896 3284 1904
rect 3276 1876 3284 1884
rect 3260 1856 3268 1864
rect 3196 1836 3204 1844
rect 3212 1836 3220 1844
rect 3340 1896 3348 1904
rect 3356 1896 3364 1904
rect 3452 2356 3460 2364
rect 3436 2316 3444 2324
rect 3484 2376 3492 2384
rect 3484 2336 3492 2344
rect 3452 2296 3460 2304
rect 3436 2256 3444 2264
rect 3404 2176 3412 2184
rect 3404 2156 3412 2164
rect 3452 2156 3460 2164
rect 3436 2136 3444 2144
rect 3532 2596 3540 2604
rect 3644 2756 3652 2764
rect 3644 2736 3652 2744
rect 3724 3696 3732 3704
rect 3756 3736 3764 3744
rect 3788 3740 3796 3744
rect 3788 3736 3796 3740
rect 3772 3696 3780 3704
rect 3772 3596 3780 3604
rect 3740 3556 3748 3564
rect 3724 3536 3732 3544
rect 3740 3496 3748 3504
rect 3756 3476 3764 3484
rect 3740 3436 3748 3444
rect 3772 3396 3780 3404
rect 3756 3376 3764 3384
rect 3708 3336 3716 3344
rect 3724 3316 3732 3324
rect 3692 3296 3700 3304
rect 3676 3276 3684 3284
rect 3724 3276 3732 3284
rect 3708 3176 3716 3184
rect 3676 3116 3684 3124
rect 3676 3036 3684 3044
rect 3692 2936 3700 2944
rect 3852 3916 3860 3924
rect 3852 3896 3860 3904
rect 3836 3876 3844 3884
rect 3852 3856 3860 3864
rect 3820 3816 3828 3824
rect 3820 3796 3828 3804
rect 3884 3996 3892 4004
rect 3916 3936 3924 3944
rect 3900 3916 3908 3924
rect 3900 3876 3908 3884
rect 3916 3856 3924 3864
rect 3900 3816 3908 3824
rect 3948 3956 3956 3964
rect 4060 4296 4068 4304
rect 4124 4296 4132 4304
rect 4220 4496 4228 4504
rect 4172 4476 4180 4484
rect 4236 4476 4244 4484
rect 4284 4456 4292 4464
rect 4188 4436 4196 4444
rect 4076 4256 4084 4264
rect 4140 4256 4148 4264
rect 4172 4256 4180 4264
rect 4060 4156 4068 4164
rect 3980 4136 3988 4144
rect 3996 4116 4004 4124
rect 3980 4076 3988 4084
rect 3980 3976 3988 3984
rect 4140 4236 4148 4244
rect 4172 4216 4180 4224
rect 4124 4156 4132 4164
rect 4108 4136 4116 4144
rect 4204 4316 4212 4324
rect 4284 4316 4292 4324
rect 4220 4296 4228 4304
rect 4716 5116 4724 5124
rect 4604 5096 4612 5104
rect 4636 5096 4644 5104
rect 4572 5076 4580 5084
rect 4588 5076 4596 5084
rect 4556 5056 4564 5064
rect 4604 5056 4612 5064
rect 4572 5036 4580 5044
rect 4764 5116 4772 5124
rect 4812 5116 4820 5124
rect 4956 5296 4964 5304
rect 4956 5256 4964 5264
rect 4924 5216 4932 5224
rect 4908 5156 4916 5164
rect 4940 5156 4948 5164
rect 4860 5076 4868 5084
rect 4844 5056 4852 5064
rect 5020 5216 5028 5224
rect 5068 5316 5076 5324
rect 5116 5316 5124 5324
rect 5244 5736 5252 5744
rect 5452 5736 5460 5744
rect 5836 5756 5844 5764
rect 5996 5756 6004 5764
rect 5916 5736 5924 5744
rect 5436 5696 5444 5704
rect 5516 5696 5524 5704
rect 5532 5696 5540 5704
rect 5612 5696 5620 5704
rect 5276 5636 5284 5644
rect 5324 5576 5332 5584
rect 5356 5576 5364 5584
rect 5228 5536 5236 5544
rect 5292 5536 5300 5544
rect 5420 5576 5428 5584
rect 5436 5576 5444 5584
rect 5404 5556 5412 5564
rect 5356 5536 5364 5544
rect 5212 5496 5220 5504
rect 5324 5496 5332 5504
rect 5164 5476 5172 5484
rect 5196 5476 5204 5484
rect 5388 5516 5396 5524
rect 5372 5496 5380 5504
rect 5916 5716 5924 5724
rect 5996 5718 6004 5724
rect 5996 5716 6004 5718
rect 5900 5696 5908 5704
rect 5596 5556 5604 5564
rect 5788 5556 5796 5564
rect 5804 5556 5812 5564
rect 5452 5536 5460 5544
rect 5484 5536 5492 5544
rect 5548 5536 5556 5544
rect 5692 5536 5700 5544
rect 5516 5516 5524 5524
rect 5468 5496 5476 5504
rect 5228 5456 5236 5464
rect 5244 5456 5252 5464
rect 5340 5456 5348 5464
rect 5356 5456 5364 5464
rect 5404 5456 5412 5464
rect 5164 5316 5172 5324
rect 5100 5296 5108 5304
rect 5132 5296 5140 5304
rect 5180 5296 5188 5304
rect 5164 5276 5172 5284
rect 5084 5256 5092 5264
rect 5132 5256 5140 5264
rect 5148 5196 5156 5204
rect 4988 5176 4996 5184
rect 5020 5156 5028 5164
rect 4892 5096 4900 5104
rect 4956 5096 4964 5104
rect 5004 5096 5012 5104
rect 4940 5076 4948 5084
rect 4732 5036 4740 5044
rect 4796 5036 4804 5044
rect 4876 5036 4884 5044
rect 5068 5076 5076 5084
rect 4988 5056 4996 5064
rect 5036 5056 5044 5064
rect 4988 5036 4996 5044
rect 5036 5036 5044 5044
rect 5084 5036 5092 5044
rect 5132 5036 5140 5044
rect 5228 5336 5236 5344
rect 5228 5316 5236 5324
rect 5596 5476 5604 5484
rect 5612 5456 5620 5464
rect 5404 5436 5412 5444
rect 5532 5436 5540 5444
rect 5564 5436 5572 5444
rect 5516 5416 5524 5424
rect 5708 5516 5716 5524
rect 5932 5576 5940 5584
rect 5932 5556 5940 5564
rect 5980 5536 5988 5544
rect 5676 5496 5684 5504
rect 5836 5496 5844 5504
rect 5788 5476 5796 5484
rect 5724 5456 5732 5464
rect 5900 5456 5908 5464
rect 5804 5416 5812 5424
rect 5612 5376 5620 5384
rect 5660 5376 5668 5384
rect 6012 5456 6020 5464
rect 5996 5376 6004 5384
rect 6060 5696 6068 5704
rect 6076 5536 6084 5544
rect 6060 5476 6068 5484
rect 5852 5356 5860 5364
rect 5948 5356 5956 5364
rect 5980 5356 5988 5364
rect 6060 5356 6068 5364
rect 5292 5336 5300 5344
rect 5340 5336 5348 5344
rect 5308 5316 5316 5324
rect 5420 5336 5428 5344
rect 5532 5336 5540 5344
rect 5548 5336 5556 5344
rect 5692 5336 5700 5344
rect 5468 5316 5476 5324
rect 5356 5296 5364 5304
rect 5244 5276 5252 5284
rect 5212 5256 5220 5264
rect 5180 5216 5188 5224
rect 5244 5156 5252 5164
rect 5340 5236 5348 5244
rect 5484 5296 5492 5304
rect 5468 5276 5476 5284
rect 5436 5256 5444 5264
rect 5612 5316 5620 5324
rect 5708 5316 5716 5324
rect 5548 5296 5556 5304
rect 5580 5296 5588 5304
rect 5532 5276 5540 5284
rect 5452 5196 5460 5204
rect 5436 5176 5444 5184
rect 5356 5136 5364 5144
rect 5212 5116 5220 5124
rect 5244 5116 5252 5124
rect 5276 5116 5284 5124
rect 5420 5116 5428 5124
rect 5212 5096 5220 5104
rect 5196 5056 5204 5064
rect 5228 5036 5236 5044
rect 4556 4976 4564 4984
rect 4620 4976 4628 4984
rect 4716 4976 4724 4984
rect 4956 4976 4964 4984
rect 4540 4956 4548 4964
rect 4540 4936 4548 4944
rect 4572 4956 4580 4964
rect 4780 4956 4788 4964
rect 4860 4956 4868 4964
rect 4924 4956 4932 4964
rect 4636 4936 4644 4944
rect 4652 4936 4660 4944
rect 4940 4936 4948 4944
rect 5100 4936 5108 4944
rect 4732 4916 4740 4924
rect 4812 4916 4820 4924
rect 4700 4896 4708 4904
rect 4780 4896 4788 4904
rect 4908 4896 4916 4904
rect 4476 4876 4484 4884
rect 4492 4876 4500 4884
rect 4524 4876 4532 4884
rect 4604 4876 4612 4884
rect 4876 4876 4884 4884
rect 4572 4836 4580 4844
rect 4638 4806 4646 4814
rect 4652 4806 4660 4814
rect 4666 4806 4674 4814
rect 4828 4796 4836 4804
rect 5020 4916 5028 4924
rect 4972 4896 4980 4904
rect 4988 4896 4996 4904
rect 4988 4796 4996 4804
rect 5052 4916 5060 4924
rect 5036 4896 5044 4904
rect 5084 4896 5092 4904
rect 5036 4856 5044 4864
rect 4796 4776 4804 4784
rect 4844 4776 4852 4784
rect 5020 4776 5028 4784
rect 4572 4756 4580 4764
rect 4604 4756 4612 4764
rect 4476 4736 4484 4744
rect 4556 4736 4564 4744
rect 4492 4716 4500 4724
rect 4460 4696 4468 4704
rect 4508 4696 4516 4704
rect 4476 4676 4484 4684
rect 4460 4656 4468 4664
rect 4444 4616 4452 4624
rect 4524 4676 4532 4684
rect 4540 4596 4548 4604
rect 4620 4736 4628 4744
rect 4636 4716 4644 4724
rect 4748 4696 4756 4704
rect 4652 4656 4660 4664
rect 4604 4596 4612 4604
rect 4780 4696 4788 4704
rect 5148 4896 5156 4904
rect 5212 4916 5220 4924
rect 5500 5256 5508 5264
rect 5612 5256 5620 5264
rect 5676 5296 5684 5304
rect 5788 5336 5796 5344
rect 5756 5316 5764 5324
rect 5820 5316 5828 5324
rect 5884 5316 5892 5324
rect 5916 5316 5924 5324
rect 5660 5276 5668 5284
rect 5740 5276 5748 5284
rect 5852 5296 5860 5304
rect 5564 5236 5572 5244
rect 5516 5196 5524 5204
rect 5484 5176 5492 5184
rect 5500 5136 5508 5144
rect 5548 5136 5556 5144
rect 5628 5236 5636 5244
rect 5740 5256 5748 5264
rect 5804 5276 5812 5284
rect 5852 5276 5860 5284
rect 5772 5256 5780 5264
rect 5676 5156 5684 5164
rect 5740 5156 5748 5164
rect 6012 5336 6020 5344
rect 6012 5316 6020 5324
rect 6044 5318 6052 5324
rect 6044 5316 6052 5318
rect 5516 5116 5524 5124
rect 5612 5116 5620 5124
rect 5708 5116 5716 5124
rect 5820 5116 5828 5124
rect 5868 5116 5876 5124
rect 5948 5116 5956 5124
rect 5340 5056 5348 5064
rect 5260 5036 5268 5044
rect 5292 5036 5300 5044
rect 5340 5036 5348 5044
rect 5260 5016 5268 5024
rect 5244 4916 5252 4924
rect 5148 4876 5156 4884
rect 5196 4796 5204 4804
rect 4988 4736 4996 4744
rect 4812 4676 4820 4684
rect 4860 4676 4868 4684
rect 4876 4676 4884 4684
rect 4764 4656 4772 4664
rect 4828 4656 4836 4664
rect 4764 4636 4772 4644
rect 5036 4696 5044 4704
rect 4972 4656 4980 4664
rect 4924 4636 4932 4644
rect 4908 4616 4916 4624
rect 4972 4616 4980 4624
rect 5116 4736 5124 4744
rect 5244 4736 5252 4744
rect 5244 4716 5252 4724
rect 5068 4696 5076 4704
rect 5052 4656 5060 4664
rect 5052 4636 5060 4644
rect 5020 4616 5028 4624
rect 4988 4596 4996 4604
rect 4492 4576 4500 4584
rect 4588 4576 4596 4584
rect 4924 4576 4932 4584
rect 4316 4536 4324 4544
rect 4396 4536 4404 4544
rect 4476 4536 4484 4544
rect 4860 4556 4868 4564
rect 5004 4556 5012 4564
rect 4716 4536 4724 4544
rect 4828 4536 4836 4544
rect 4908 4536 4916 4544
rect 5020 4536 5028 4544
rect 4540 4516 4548 4524
rect 4348 4456 4356 4464
rect 4508 4456 4516 4464
rect 4524 4436 4532 4444
rect 4412 4416 4420 4424
rect 4380 4316 4388 4324
rect 4364 4296 4372 4304
rect 4220 4136 4228 4144
rect 4204 4116 4212 4124
rect 4108 4096 4116 4104
rect 4140 4096 4148 4104
rect 4172 4096 4180 4104
rect 4076 4056 4084 4064
rect 4140 4076 4148 4084
rect 4124 4056 4132 4064
rect 4124 3996 4132 4004
rect 4092 3976 4100 3984
rect 4012 3956 4020 3964
rect 4044 3956 4052 3964
rect 4060 3956 4068 3964
rect 4284 4136 4292 4144
rect 4252 4096 4260 4104
rect 4188 3936 4196 3944
rect 4252 3936 4260 3944
rect 4044 3916 4052 3924
rect 4076 3916 4084 3924
rect 4156 3916 4164 3924
rect 4172 3916 4180 3924
rect 4220 3916 4228 3924
rect 3980 3896 3988 3904
rect 4060 3896 4068 3904
rect 4092 3896 4100 3904
rect 4108 3896 4116 3904
rect 4044 3876 4052 3884
rect 3964 3816 3972 3824
rect 4236 3896 4244 3904
rect 4268 3896 4276 3904
rect 4156 3816 4164 3824
rect 4188 3816 4196 3824
rect 4332 4116 4340 4124
rect 4348 4096 4356 4104
rect 4380 4136 4388 4144
rect 4572 4516 4580 4524
rect 4716 4516 4724 4524
rect 4796 4516 4804 4524
rect 4620 4496 4628 4504
rect 4700 4496 4708 4504
rect 4764 4496 4772 4504
rect 4556 4456 4564 4464
rect 4540 4416 4548 4424
rect 4638 4406 4646 4414
rect 4652 4406 4660 4414
rect 4666 4406 4674 4414
rect 4764 4476 4772 4484
rect 4444 4316 4452 4324
rect 4428 4276 4436 4284
rect 4684 4296 4692 4304
rect 4492 4276 4500 4284
rect 4460 4256 4468 4264
rect 4588 4256 4596 4264
rect 4604 4256 4612 4264
rect 4556 4236 4564 4244
rect 4732 4196 4740 4204
rect 4572 4176 4580 4184
rect 4604 4176 4612 4184
rect 4460 4156 4468 4164
rect 4412 4116 4420 4124
rect 4444 4116 4452 4124
rect 4428 4096 4436 4104
rect 4316 4076 4324 4084
rect 4396 4076 4404 4084
rect 4396 4036 4404 4044
rect 4316 3976 4324 3984
rect 4300 3956 4308 3964
rect 4364 3956 4372 3964
rect 4332 3936 4340 3944
rect 4348 3916 4356 3924
rect 4316 3896 4324 3904
rect 4332 3896 4340 3904
rect 4444 3956 4452 3964
rect 4524 4156 4532 4164
rect 4556 4156 4564 4164
rect 4476 4076 4484 4084
rect 4428 3936 4436 3944
rect 4460 3916 4468 3924
rect 4396 3896 4404 3904
rect 4316 3876 4324 3884
rect 4332 3876 4340 3884
rect 4284 3856 4292 3864
rect 4236 3776 4244 3784
rect 4284 3776 4292 3784
rect 4076 3756 4084 3764
rect 4156 3756 4164 3764
rect 3948 3736 3956 3744
rect 4012 3736 4020 3744
rect 3836 3636 3844 3644
rect 3836 3596 3844 3604
rect 4220 3736 4228 3744
rect 4252 3736 4260 3744
rect 3996 3716 4004 3724
rect 4076 3716 4084 3724
rect 4108 3716 4116 3724
rect 3964 3576 3972 3584
rect 3932 3556 3940 3564
rect 3868 3496 3876 3504
rect 3852 3456 3860 3464
rect 3868 3436 3876 3444
rect 3836 3416 3844 3424
rect 3820 3396 3828 3404
rect 3964 3456 3972 3464
rect 4044 3696 4052 3704
rect 4076 3696 4084 3704
rect 4156 3696 4164 3704
rect 4092 3676 4100 3684
rect 4140 3676 4148 3684
rect 4204 3676 4212 3684
rect 4188 3656 4196 3664
rect 4236 3656 4244 3664
rect 4204 3636 4212 3644
rect 4300 3696 4308 3704
rect 4060 3556 4068 3564
rect 4172 3556 4180 3564
rect 4300 3536 4308 3544
rect 4076 3516 4084 3524
rect 4156 3516 4164 3524
rect 4268 3516 4276 3524
rect 4204 3496 4212 3504
rect 4156 3476 4164 3484
rect 4108 3456 4116 3464
rect 4012 3436 4020 3444
rect 4124 3436 4132 3444
rect 3996 3416 4004 3424
rect 3900 3396 3908 3404
rect 4044 3396 4052 3404
rect 4204 3396 4212 3404
rect 3852 3376 3860 3384
rect 4220 3376 4228 3384
rect 4220 3356 4228 3364
rect 3740 3196 3748 3204
rect 3772 3196 3780 3204
rect 3756 3156 3764 3164
rect 3932 3316 3940 3324
rect 3996 3316 4004 3324
rect 3980 3296 3988 3304
rect 3964 3236 3972 3244
rect 3916 3216 3924 3224
rect 3900 3196 3908 3204
rect 3820 3176 3828 3184
rect 3868 3176 3876 3184
rect 3852 3156 3860 3164
rect 3916 3176 3924 3184
rect 4108 3336 4116 3344
rect 4252 3436 4260 3444
rect 4060 3316 4068 3324
rect 4108 3316 4116 3324
rect 4236 3316 4244 3324
rect 4028 3296 4036 3304
rect 4012 3236 4020 3244
rect 4060 3216 4068 3224
rect 3948 3156 3956 3164
rect 4028 3136 4036 3144
rect 3868 3116 3876 3124
rect 3884 3116 3892 3124
rect 4012 3116 4020 3124
rect 4076 3196 4084 3204
rect 3900 3096 3908 3104
rect 3996 3096 4004 3104
rect 4028 3096 4036 3104
rect 3756 3076 3764 3084
rect 3788 3076 3796 3084
rect 3836 3076 3844 3084
rect 3852 3076 3860 3084
rect 3900 3076 3908 3084
rect 3740 3036 3748 3044
rect 3724 2896 3732 2904
rect 3676 2856 3684 2864
rect 3724 2776 3732 2784
rect 3660 2716 3668 2724
rect 3612 2656 3620 2664
rect 3628 2656 3636 2664
rect 3612 2616 3620 2624
rect 3612 2576 3620 2584
rect 3532 2536 3540 2544
rect 3596 2536 3604 2544
rect 3548 2496 3556 2504
rect 3532 2476 3540 2484
rect 3516 2416 3524 2424
rect 3516 2316 3524 2324
rect 3532 2316 3540 2324
rect 3500 2296 3508 2304
rect 3484 2276 3492 2284
rect 3580 2476 3588 2484
rect 3644 2556 3652 2564
rect 3628 2536 3636 2544
rect 3612 2456 3620 2464
rect 3580 2416 3588 2424
rect 3612 2376 3620 2384
rect 3612 2336 3620 2344
rect 3596 2316 3604 2324
rect 3740 2756 3748 2764
rect 3708 2616 3716 2624
rect 3772 3056 3780 3064
rect 3868 3036 3876 3044
rect 3916 3036 3924 3044
rect 3852 2996 3860 3004
rect 3788 2976 3796 2984
rect 3836 2936 3844 2944
rect 3868 2936 3876 2944
rect 3820 2916 3828 2924
rect 3836 2896 3844 2904
rect 3804 2856 3812 2864
rect 3772 2756 3780 2764
rect 3868 2856 3876 2864
rect 3836 2836 3844 2844
rect 3884 2836 3892 2844
rect 3804 2736 3812 2744
rect 3820 2736 3828 2744
rect 3772 2716 3780 2724
rect 3772 2696 3780 2704
rect 3820 2696 3828 2704
rect 4092 3116 4100 3124
rect 4092 3096 4100 3104
rect 4092 3076 4100 3084
rect 3964 3056 3972 3064
rect 4044 3036 4052 3044
rect 3948 3016 3956 3024
rect 4156 3156 4164 3164
rect 4172 3136 4180 3144
rect 4236 3196 4244 3204
rect 4204 3156 4212 3164
rect 4156 3116 4164 3124
rect 4124 3096 4132 3104
rect 4108 3056 4116 3064
rect 4140 3016 4148 3024
rect 4124 2996 4132 3004
rect 4012 2976 4020 2984
rect 3948 2936 3956 2944
rect 4028 2956 4036 2964
rect 4092 2956 4100 2964
rect 4044 2936 4052 2944
rect 3980 2896 3988 2904
rect 4012 2876 4020 2884
rect 3932 2856 3940 2864
rect 3948 2776 3956 2784
rect 3996 2776 4004 2784
rect 3932 2716 3940 2724
rect 3964 2716 3972 2724
rect 3884 2696 3892 2704
rect 3916 2696 3924 2704
rect 3836 2676 3844 2684
rect 3916 2676 3924 2684
rect 3836 2656 3844 2664
rect 3756 2616 3764 2624
rect 3820 2616 3828 2624
rect 3740 2576 3748 2584
rect 3724 2556 3732 2564
rect 3708 2536 3716 2544
rect 3740 2536 3748 2544
rect 3676 2496 3684 2504
rect 3660 2456 3668 2464
rect 3644 2336 3652 2344
rect 3596 2276 3604 2284
rect 3628 2276 3636 2284
rect 3484 2256 3492 2264
rect 3548 2256 3556 2264
rect 3420 2116 3428 2124
rect 3468 2076 3476 2084
rect 3436 2056 3444 2064
rect 3388 1916 3396 1924
rect 3324 1876 3332 1884
rect 3372 1876 3380 1884
rect 3308 1856 3316 1864
rect 3228 1776 3236 1784
rect 3276 1776 3284 1784
rect 3196 1756 3204 1764
rect 3212 1756 3220 1764
rect 3276 1756 3284 1764
rect 3292 1756 3300 1764
rect 3260 1736 3268 1744
rect 3276 1736 3284 1744
rect 3228 1696 3236 1704
rect 3292 1696 3300 1704
rect 3196 1636 3204 1644
rect 3228 1616 3236 1624
rect 3276 1616 3284 1624
rect 3132 1556 3140 1564
rect 3020 1476 3028 1484
rect 3036 1476 3044 1484
rect 2988 1456 2996 1464
rect 3004 1456 3012 1464
rect 2924 1416 2932 1424
rect 2908 1336 2916 1344
rect 2908 1316 2916 1324
rect 2892 1296 2900 1304
rect 2844 1236 2852 1244
rect 2812 1196 2820 1204
rect 2828 1196 2836 1204
rect 2764 1136 2772 1144
rect 2620 1096 2628 1104
rect 2684 1096 2692 1104
rect 2732 1096 2740 1104
rect 2780 1116 2788 1124
rect 2972 1396 2980 1404
rect 2956 1376 2964 1384
rect 2972 1336 2980 1344
rect 3004 1416 3012 1424
rect 3132 1476 3140 1484
rect 3148 1476 3156 1484
rect 3196 1496 3204 1504
rect 3244 1576 3252 1584
rect 3260 1556 3268 1564
rect 3244 1536 3252 1544
rect 3260 1496 3268 1504
rect 3180 1476 3188 1484
rect 3164 1456 3172 1464
rect 3084 1416 3092 1424
rect 3118 1406 3126 1414
rect 3132 1406 3140 1414
rect 3146 1406 3154 1414
rect 3196 1436 3204 1444
rect 3212 1436 3220 1444
rect 3180 1396 3188 1404
rect 3036 1376 3044 1384
rect 3068 1336 3076 1344
rect 3084 1316 3092 1324
rect 3180 1316 3188 1324
rect 3228 1316 3236 1324
rect 3308 1556 3316 1564
rect 3340 1816 3348 1824
rect 3356 1796 3364 1804
rect 3340 1736 3348 1744
rect 3452 1836 3460 1844
rect 3452 1776 3460 1784
rect 3388 1756 3396 1764
rect 3388 1736 3396 1744
rect 3372 1696 3380 1704
rect 3404 1676 3412 1684
rect 3388 1576 3396 1584
rect 3372 1556 3380 1564
rect 3340 1536 3348 1544
rect 3388 1476 3396 1484
rect 3340 1436 3348 1444
rect 3452 1656 3460 1664
rect 3452 1576 3460 1584
rect 3516 2176 3524 2184
rect 3532 2176 3540 2184
rect 3500 2076 3508 2084
rect 3484 1956 3492 1964
rect 3500 1956 3508 1964
rect 3516 1916 3524 1924
rect 3612 2256 3620 2264
rect 3564 2176 3572 2184
rect 3612 2176 3620 2184
rect 3564 2156 3572 2164
rect 3596 2156 3604 2164
rect 3500 1896 3508 1904
rect 3548 1896 3556 1904
rect 3484 1856 3492 1864
rect 3548 1856 3556 1864
rect 3420 1516 3428 1524
rect 3436 1476 3444 1484
rect 3324 1416 3332 1424
rect 3404 1416 3412 1424
rect 3372 1396 3380 1404
rect 3356 1376 3364 1384
rect 3020 1296 3028 1304
rect 3212 1296 3220 1304
rect 3244 1296 3252 1304
rect 2940 1236 2948 1244
rect 2924 1216 2932 1224
rect 2860 1156 2868 1164
rect 2876 1156 2884 1164
rect 3020 1156 3028 1164
rect 2908 1136 2916 1144
rect 2924 1136 2932 1144
rect 2892 1116 2900 1124
rect 2924 1116 2932 1124
rect 2972 1116 2980 1124
rect 3020 1116 3028 1124
rect 3340 1296 3348 1304
rect 3276 1256 3284 1264
rect 3292 1256 3300 1264
rect 3164 1236 3172 1244
rect 3084 1176 3092 1184
rect 3052 1156 3060 1164
rect 2796 1096 2804 1104
rect 2812 1096 2820 1104
rect 2892 1096 2900 1104
rect 2908 1096 2916 1104
rect 2988 1096 2996 1104
rect 3036 1096 3044 1104
rect 2956 1036 2964 1044
rect 3036 1036 3044 1044
rect 2732 1016 2740 1024
rect 2908 1016 2916 1024
rect 2588 996 2596 1004
rect 2620 976 2628 984
rect 2636 936 2644 944
rect 2588 896 2596 904
rect 2652 896 2660 904
rect 2588 876 2596 884
rect 2652 876 2660 884
rect 2684 856 2692 864
rect 2572 836 2580 844
rect 2540 736 2548 744
rect 2508 716 2516 724
rect 2524 716 2532 724
rect 2332 696 2340 704
rect 2364 676 2372 684
rect 2332 656 2340 664
rect 2412 656 2420 664
rect 2316 616 2324 624
rect 2380 616 2388 624
rect 2348 596 2356 604
rect 2476 656 2484 664
rect 2460 636 2468 644
rect 2508 636 2516 644
rect 2524 636 2532 644
rect 2396 556 2404 564
rect 2428 556 2436 564
rect 2444 556 2452 564
rect 2508 556 2516 564
rect 2540 556 2548 564
rect 2556 556 2564 564
rect 2268 536 2276 544
rect 2220 516 2228 524
rect 2156 496 2164 504
rect 2220 496 2228 504
rect 2236 496 2244 504
rect 2284 496 2292 504
rect 2076 376 2084 384
rect 2124 376 2132 384
rect 1884 356 1892 364
rect 1948 356 1956 364
rect 1836 336 1844 344
rect 1820 296 1828 304
rect 1900 296 1908 304
rect 1820 216 1828 224
rect 1852 276 1860 284
rect 2396 516 2404 524
rect 2268 476 2276 484
rect 2380 476 2388 484
rect 2300 436 2308 444
rect 2236 336 2244 344
rect 2060 316 2068 324
rect 2252 316 2260 324
rect 2076 276 2084 284
rect 1932 256 1940 264
rect 1852 236 1860 244
rect 1852 216 1860 224
rect 1836 176 1844 184
rect 1852 156 1860 164
rect 1532 136 1540 144
rect 1628 136 1636 144
rect 1516 116 1524 124
rect 1452 96 1460 104
rect 1484 96 1492 104
rect 1566 6 1574 14
rect 1580 6 1588 14
rect 1594 6 1602 14
rect 1916 156 1924 164
rect 1948 156 1956 164
rect 1980 156 1988 164
rect 2028 156 2036 164
rect 2044 156 2052 164
rect 2076 156 2084 164
rect 1916 136 1924 144
rect 1884 116 1892 124
rect 1932 96 1940 104
rect 1948 96 1956 104
rect 1964 96 1972 104
rect 2012 116 2020 124
rect 2044 116 2052 124
rect 1996 96 2004 104
rect 2108 216 2116 224
rect 2188 276 2196 284
rect 2284 276 2292 284
rect 2156 256 2164 264
rect 2188 256 2196 264
rect 2236 256 2244 264
rect 2140 196 2148 204
rect 2348 396 2356 404
rect 2332 256 2340 264
rect 2524 536 2532 544
rect 2508 516 2516 524
rect 2700 816 2708 824
rect 2668 756 2676 764
rect 2716 756 2724 764
rect 2604 656 2612 664
rect 2700 736 2708 744
rect 2668 656 2676 664
rect 2652 636 2660 644
rect 2684 616 2692 624
rect 2668 596 2676 604
rect 2988 996 2996 1004
rect 3020 996 3028 1004
rect 2860 976 2868 984
rect 2828 956 2836 964
rect 3036 956 3044 964
rect 2860 916 2868 924
rect 2860 896 2868 904
rect 2908 896 2916 904
rect 2796 876 2804 884
rect 2748 856 2756 864
rect 2780 856 2788 864
rect 2748 796 2756 804
rect 2796 796 2804 804
rect 2764 776 2772 784
rect 2796 756 2804 764
rect 3100 1116 3108 1124
rect 3292 1196 3300 1204
rect 3324 1196 3332 1204
rect 3228 1176 3236 1184
rect 3308 1176 3316 1184
rect 3196 1156 3204 1164
rect 3420 1396 3428 1404
rect 3420 1376 3428 1384
rect 3468 1516 3476 1524
rect 3516 1836 3524 1844
rect 3500 1776 3508 1784
rect 3596 2076 3604 2084
rect 3580 2036 3588 2044
rect 3660 2196 3668 2204
rect 3676 2136 3684 2144
rect 3644 2096 3652 2104
rect 3676 2076 3684 2084
rect 3628 2056 3636 2064
rect 3676 2056 3684 2064
rect 3612 1956 3620 1964
rect 3676 1956 3684 1964
rect 3580 1916 3588 1924
rect 3644 1896 3652 1904
rect 3660 1896 3668 1904
rect 3580 1856 3588 1864
rect 3612 1796 3620 1804
rect 3596 1776 3604 1784
rect 3564 1756 3572 1764
rect 3548 1696 3556 1704
rect 3532 1616 3540 1624
rect 3548 1616 3556 1624
rect 3580 1536 3588 1544
rect 3644 1796 3652 1804
rect 3660 1776 3668 1784
rect 3612 1756 3620 1764
rect 3628 1756 3636 1764
rect 3644 1756 3652 1764
rect 3612 1656 3620 1664
rect 3644 1636 3652 1644
rect 3596 1476 3604 1484
rect 3580 1436 3588 1444
rect 3516 1416 3524 1424
rect 3532 1416 3540 1424
rect 3500 1376 3508 1384
rect 3452 1356 3460 1364
rect 3452 1336 3460 1344
rect 3484 1336 3492 1344
rect 3420 1316 3428 1324
rect 3532 1336 3540 1344
rect 3468 1256 3476 1264
rect 3500 1276 3508 1284
rect 3516 1276 3524 1284
rect 3372 1216 3380 1224
rect 3244 1136 3252 1144
rect 3340 1136 3348 1144
rect 3356 1136 3364 1144
rect 3212 1116 3220 1124
rect 3404 1136 3412 1144
rect 3260 1116 3268 1124
rect 3308 1116 3316 1124
rect 3324 1116 3332 1124
rect 3468 1116 3476 1124
rect 3532 1216 3540 1224
rect 3516 1176 3524 1184
rect 3580 1376 3588 1384
rect 3756 2516 3764 2524
rect 3708 2496 3716 2504
rect 3724 2496 3732 2504
rect 3724 2456 3732 2464
rect 3740 2456 3748 2464
rect 3724 2416 3732 2424
rect 3724 2296 3732 2304
rect 3724 2276 3732 2284
rect 3788 2516 3796 2524
rect 4092 2916 4100 2924
rect 4060 2856 4068 2864
rect 4076 2736 4084 2744
rect 4092 2736 4100 2744
rect 4124 2736 4132 2744
rect 4012 2716 4020 2724
rect 4028 2716 4036 2724
rect 4060 2716 4068 2724
rect 3980 2696 3988 2704
rect 4044 2696 4052 2704
rect 3948 2676 3956 2684
rect 3964 2656 3972 2664
rect 4108 2716 4116 2724
rect 4092 2696 4100 2704
rect 4028 2656 4036 2664
rect 4108 2656 4116 2664
rect 4044 2636 4052 2644
rect 4092 2636 4100 2644
rect 3980 2576 3988 2584
rect 3884 2556 3892 2564
rect 3932 2556 3940 2564
rect 3836 2536 3844 2544
rect 3964 2536 3972 2544
rect 3996 2536 4004 2544
rect 3900 2516 3908 2524
rect 3916 2516 3924 2524
rect 3820 2476 3828 2484
rect 3884 2476 3892 2484
rect 3804 2456 3812 2464
rect 3820 2456 3828 2464
rect 3868 2456 3876 2464
rect 3772 2436 3780 2444
rect 3980 2436 3988 2444
rect 4012 2516 4020 2524
rect 4060 2576 4068 2584
rect 4060 2536 4068 2544
rect 4076 2496 4084 2504
rect 3996 2396 4004 2404
rect 3836 2376 3844 2384
rect 3756 2336 3764 2344
rect 3772 2336 3780 2344
rect 3820 2336 3828 2344
rect 3884 2316 3892 2324
rect 3900 2316 3908 2324
rect 3964 2316 3972 2324
rect 3740 2236 3748 2244
rect 3756 2236 3764 2244
rect 3916 2296 3924 2304
rect 4044 2396 4052 2404
rect 4060 2316 4068 2324
rect 3964 2276 3972 2284
rect 3916 2256 3924 2264
rect 4012 2276 4020 2284
rect 3836 2236 3844 2244
rect 3996 2236 4004 2244
rect 4092 2256 4100 2264
rect 3788 2216 3796 2224
rect 4028 2216 4036 2224
rect 4172 3096 4180 3104
rect 4300 3496 4308 3504
rect 4396 3816 4404 3824
rect 4428 3816 4436 3824
rect 4396 3796 4404 3804
rect 4508 3896 4516 3904
rect 4524 3816 4532 3824
rect 4876 4516 4884 4524
rect 5228 4676 5236 4684
rect 5116 4636 5124 4644
rect 5212 4616 5220 4624
rect 5100 4596 5108 4604
rect 5084 4576 5092 4584
rect 5116 4576 5124 4584
rect 5164 4576 5172 4584
rect 5132 4536 5140 4544
rect 5244 4536 5252 4544
rect 5132 4516 5140 4524
rect 5228 4516 5236 4524
rect 4860 4496 4868 4504
rect 5100 4496 5108 4504
rect 4844 4316 4852 4324
rect 4844 4256 4852 4264
rect 4972 4476 4980 4484
rect 5052 4336 5060 4344
rect 5084 4336 5092 4344
rect 5244 4336 5252 4344
rect 4876 4316 4884 4324
rect 5132 4316 5140 4324
rect 5244 4316 5252 4324
rect 4924 4276 4932 4284
rect 4892 4256 4900 4264
rect 4876 4236 4884 4244
rect 4844 4176 4852 4184
rect 4828 4156 4836 4164
rect 4604 4096 4612 4104
rect 4780 4136 4788 4144
rect 4940 4256 4948 4264
rect 5116 4296 5124 4304
rect 4988 4276 4996 4284
rect 4956 4236 4964 4244
rect 5004 4156 5012 4164
rect 4956 4136 4964 4144
rect 4908 4116 4916 4124
rect 4924 4116 4932 4124
rect 4764 4096 4772 4104
rect 4620 4076 4628 4084
rect 4668 4076 4676 4084
rect 4700 4076 4708 4084
rect 4638 4006 4646 4014
rect 4652 4006 4660 4014
rect 4666 4006 4674 4014
rect 4588 3976 4596 3984
rect 4844 4076 4852 4084
rect 4780 4036 4788 4044
rect 4780 3976 4788 3984
rect 4940 4096 4948 4104
rect 4988 4096 4996 4104
rect 4956 4076 4964 4084
rect 4908 4056 4916 4064
rect 5228 4276 5236 4284
rect 5132 4256 5140 4264
rect 5100 4176 5108 4184
rect 5036 4136 5044 4144
rect 5100 4136 5108 4144
rect 5036 4116 5044 4124
rect 5052 4116 5060 4124
rect 5020 4056 5028 4064
rect 4972 4036 4980 4044
rect 5004 4036 5012 4044
rect 5004 4016 5012 4024
rect 5052 4056 5060 4064
rect 5116 4056 5124 4064
rect 5100 4016 5108 4024
rect 5244 4216 5252 4224
rect 5164 4196 5172 4204
rect 5228 4196 5236 4204
rect 5164 4176 5172 4184
rect 5148 4156 5156 4164
rect 5244 4156 5252 4164
rect 5180 4136 5188 4144
rect 5164 4116 5172 4124
rect 5244 4116 5252 4124
rect 4892 3976 4900 3984
rect 5244 4096 5252 4104
rect 5324 4956 5332 4964
rect 5356 4956 5364 4964
rect 5292 4916 5300 4924
rect 5276 4896 5284 4904
rect 5308 4716 5316 4724
rect 5292 4676 5300 4684
rect 5388 4916 5396 4924
rect 5372 4896 5380 4904
rect 5532 5096 5540 5104
rect 5548 5076 5556 5084
rect 5580 5080 5588 5084
rect 5580 5076 5588 5080
rect 5660 5096 5668 5104
rect 5724 5096 5732 5104
rect 5900 5096 5908 5104
rect 5804 5076 5812 5084
rect 5836 5076 5844 5084
rect 5580 4956 5588 4964
rect 5420 4936 5428 4944
rect 5500 4936 5508 4944
rect 5548 4936 5556 4944
rect 5580 4936 5588 4944
rect 5436 4916 5444 4924
rect 5340 4876 5348 4884
rect 5292 4656 5300 4664
rect 5324 4656 5332 4664
rect 5276 4496 5284 4504
rect 5356 4676 5364 4684
rect 5356 4656 5364 4664
rect 5356 4616 5364 4624
rect 5308 4540 5316 4544
rect 5308 4536 5316 4540
rect 5372 4556 5380 4564
rect 5372 4516 5380 4524
rect 5404 4856 5412 4864
rect 5468 4876 5476 4884
rect 5452 4856 5460 4864
rect 5436 4836 5444 4844
rect 5436 4816 5444 4824
rect 5516 4736 5524 4744
rect 5484 4716 5492 4724
rect 5420 4696 5428 4704
rect 5468 4696 5476 4704
rect 5500 4696 5508 4704
rect 5532 4716 5540 4724
rect 5596 4816 5604 4824
rect 5740 4956 5748 4964
rect 5788 4956 5796 4964
rect 5644 4736 5652 4744
rect 5692 4896 5700 4904
rect 5740 4896 5748 4904
rect 5804 4916 5812 4924
rect 5660 4716 5668 4724
rect 5708 4696 5716 4704
rect 5564 4676 5572 4684
rect 5580 4676 5588 4684
rect 5692 4676 5700 4684
rect 5484 4656 5492 4664
rect 5580 4656 5588 4664
rect 5436 4636 5444 4644
rect 5596 4616 5604 4624
rect 5484 4576 5492 4584
rect 5404 4536 5412 4544
rect 5452 4536 5460 4544
rect 5436 4336 5444 4344
rect 5276 4316 5284 4324
rect 5292 4296 5300 4304
rect 5276 4276 5284 4284
rect 5276 4236 5284 4244
rect 5260 4056 5268 4064
rect 5084 3956 5092 3964
rect 5196 3956 5204 3964
rect 4700 3916 4708 3924
rect 4716 3916 4724 3924
rect 4828 3916 4836 3924
rect 4588 3896 4596 3904
rect 4828 3876 4836 3884
rect 4860 3876 4868 3884
rect 4892 3876 4900 3884
rect 4588 3856 4596 3864
rect 4540 3796 4548 3804
rect 4556 3796 4564 3804
rect 4492 3776 4500 3784
rect 4476 3756 4484 3764
rect 4508 3756 4516 3764
rect 4604 3836 4612 3844
rect 4604 3796 4612 3804
rect 4652 3816 4660 3824
rect 4732 3836 4740 3844
rect 4780 3796 4788 3804
rect 4700 3776 4708 3784
rect 4716 3776 4724 3784
rect 4332 3716 4340 3724
rect 4412 3716 4420 3724
rect 4332 3696 4340 3704
rect 4396 3696 4404 3704
rect 4364 3636 4372 3644
rect 4332 3576 4340 3584
rect 4364 3556 4372 3564
rect 4444 3556 4452 3564
rect 4412 3536 4420 3544
rect 4476 3536 4484 3544
rect 4636 3756 4644 3764
rect 4636 3656 4644 3664
rect 4716 3716 4724 3724
rect 4796 3776 4804 3784
rect 4748 3656 4756 3664
rect 4700 3616 4708 3624
rect 4638 3606 4646 3614
rect 4652 3606 4660 3614
rect 4666 3606 4674 3614
rect 4588 3576 4596 3584
rect 4684 3576 4692 3584
rect 4572 3556 4580 3564
rect 4540 3536 4548 3544
rect 4492 3496 4500 3504
rect 4396 3476 4404 3484
rect 4460 3476 4468 3484
rect 4508 3476 4516 3484
rect 4540 3476 4548 3484
rect 4572 3476 4580 3484
rect 4348 3456 4356 3464
rect 4380 3456 4388 3464
rect 4460 3416 4468 3424
rect 4412 3396 4420 3404
rect 4284 3376 4292 3384
rect 4268 3356 4276 3364
rect 4268 3336 4276 3344
rect 4396 3336 4404 3344
rect 4380 3256 4388 3264
rect 4252 3116 4260 3124
rect 4764 3516 4772 3524
rect 4764 3476 4772 3484
rect 4556 3396 4564 3404
rect 4620 3396 4628 3404
rect 4604 3336 4612 3344
rect 4492 3316 4500 3324
rect 4428 3276 4436 3284
rect 4556 3316 4564 3324
rect 4588 3276 4596 3284
rect 4684 3276 4692 3284
rect 4556 3176 4564 3184
rect 4540 3156 4548 3164
rect 4540 3136 4548 3144
rect 4428 3116 4436 3124
rect 4220 3096 4228 3104
rect 4476 3096 4484 3104
rect 4188 3056 4196 3064
rect 4252 3056 4260 3064
rect 4284 3056 4292 3064
rect 4380 3056 4388 3064
rect 4348 3036 4356 3044
rect 4252 2996 4260 3004
rect 4300 2996 4308 3004
rect 4236 2936 4244 2944
rect 4348 2936 4356 2944
rect 4204 2916 4212 2924
rect 4220 2896 4228 2904
rect 4268 2876 4276 2884
rect 4188 2856 4196 2864
rect 4236 2776 4244 2784
rect 4220 2736 4228 2744
rect 4638 3206 4646 3214
rect 4652 3206 4660 3214
rect 4666 3206 4674 3214
rect 4620 3156 4628 3164
rect 4812 3736 4820 3744
rect 4844 3816 4852 3824
rect 4956 3856 4964 3864
rect 5004 3896 5012 3904
rect 5004 3876 5012 3884
rect 5212 3916 5220 3924
rect 5244 3916 5252 3924
rect 5084 3896 5092 3904
rect 5100 3896 5108 3904
rect 5148 3896 5156 3904
rect 5164 3896 5172 3904
rect 5196 3896 5204 3904
rect 5020 3856 5028 3864
rect 5068 3856 5076 3864
rect 4892 3756 4900 3764
rect 4860 3736 4868 3744
rect 4908 3736 4916 3744
rect 4940 3736 4948 3744
rect 4956 3716 4964 3724
rect 4908 3636 4916 3644
rect 4828 3596 4836 3604
rect 4828 3556 4836 3564
rect 4812 3536 4820 3544
rect 4924 3516 4932 3524
rect 4812 3476 4820 3484
rect 4844 3476 4852 3484
rect 4844 3416 4852 3424
rect 4860 3376 4868 3384
rect 4716 3356 4724 3364
rect 4828 3356 4836 3364
rect 4876 3356 4884 3364
rect 4732 3336 4740 3344
rect 4860 3336 4868 3344
rect 4716 3176 4724 3184
rect 4604 3136 4612 3144
rect 4572 3096 4580 3104
rect 4492 3076 4500 3084
rect 4524 3076 4532 3084
rect 4476 2976 4484 2984
rect 4476 2956 4484 2964
rect 4412 2936 4420 2944
rect 4300 2896 4308 2904
rect 4412 2876 4420 2884
rect 4460 2916 4468 2924
rect 4508 2936 4516 2944
rect 4492 2916 4500 2924
rect 4428 2836 4436 2844
rect 4380 2816 4388 2824
rect 4300 2776 4308 2784
rect 4332 2776 4340 2784
rect 4428 2776 4436 2784
rect 4444 2776 4452 2784
rect 4316 2756 4324 2764
rect 4284 2736 4292 2744
rect 4300 2736 4308 2744
rect 4236 2716 4244 2724
rect 4172 2696 4180 2704
rect 4300 2716 4308 2724
rect 4476 2856 4484 2864
rect 4476 2836 4484 2844
rect 4460 2756 4468 2764
rect 4572 3056 4580 3064
rect 4588 3036 4596 3044
rect 4700 3076 4708 3084
rect 4636 3056 4644 3064
rect 4620 3016 4628 3024
rect 4684 2976 4692 2984
rect 4620 2956 4628 2964
rect 4748 3116 4756 3124
rect 4844 3316 4852 3324
rect 4844 3096 4852 3104
rect 4860 3096 4868 3104
rect 4732 3076 4740 3084
rect 4780 3076 4788 3084
rect 4796 3076 4804 3084
rect 4716 3016 4724 3024
rect 4748 3056 4756 3064
rect 4748 2996 4756 3004
rect 4780 2976 4788 2984
rect 4700 2956 4708 2964
rect 4780 2956 4788 2964
rect 4540 2936 4548 2944
rect 4764 2936 4772 2944
rect 4556 2916 4564 2924
rect 4828 3056 4836 3064
rect 4796 2916 4804 2924
rect 4924 3496 4932 3504
rect 4988 3496 4996 3504
rect 4988 3476 4996 3484
rect 4908 3416 4916 3424
rect 5052 3836 5060 3844
rect 5132 3876 5140 3884
rect 5100 3856 5108 3864
rect 5132 3836 5140 3844
rect 5244 3836 5252 3844
rect 5308 4256 5316 4264
rect 5308 4156 5316 4164
rect 5324 4116 5332 4124
rect 5292 4016 5300 4024
rect 5324 3896 5332 3904
rect 5404 4216 5412 4224
rect 5420 4176 5428 4184
rect 5404 4156 5412 4164
rect 5356 4136 5364 4144
rect 5420 4096 5428 4104
rect 5356 4076 5364 4084
rect 5388 4076 5396 4084
rect 5452 4276 5460 4284
rect 5452 4116 5460 4124
rect 5404 4056 5412 4064
rect 5436 4056 5444 4064
rect 5372 3916 5380 3924
rect 5292 3836 5300 3844
rect 5388 3876 5396 3884
rect 5564 4556 5572 4564
rect 5564 4516 5572 4524
rect 5532 4396 5540 4404
rect 5548 4276 5556 4284
rect 5532 4236 5540 4244
rect 5948 5096 5956 5104
rect 5932 4956 5940 4964
rect 5836 4916 5844 4924
rect 5900 4916 5908 4924
rect 5932 4916 5940 4924
rect 5884 4896 5892 4904
rect 5820 4876 5828 4884
rect 5852 4876 5860 4884
rect 5772 4816 5780 4824
rect 5740 4776 5748 4784
rect 5772 4756 5780 4764
rect 5756 4736 5764 4744
rect 5868 4836 5876 4844
rect 5804 4756 5812 4764
rect 5852 4756 5860 4764
rect 5820 4736 5828 4744
rect 5836 4736 5844 4744
rect 5788 4716 5796 4724
rect 5772 4696 5780 4704
rect 5756 4676 5764 4684
rect 5692 4656 5700 4664
rect 5724 4656 5732 4664
rect 5740 4656 5748 4664
rect 5676 4616 5684 4624
rect 5708 4616 5716 4624
rect 5676 4556 5684 4564
rect 5788 4596 5796 4604
rect 5612 4536 5620 4544
rect 5596 4496 5604 4504
rect 5580 4356 5588 4364
rect 5612 4336 5620 4344
rect 5596 4316 5604 4324
rect 5580 4276 5588 4284
rect 5484 4076 5492 4084
rect 5484 4056 5492 4064
rect 5500 3936 5508 3944
rect 5516 3916 5524 3924
rect 5532 3876 5540 3884
rect 5580 4236 5588 4244
rect 5628 4296 5636 4304
rect 5676 4296 5684 4304
rect 5612 4276 5620 4284
rect 5660 4276 5668 4284
rect 5724 4536 5732 4544
rect 5756 4536 5764 4544
rect 5724 4496 5732 4504
rect 5708 4436 5716 4444
rect 5628 4236 5636 4244
rect 5660 4236 5668 4244
rect 5596 4216 5604 4224
rect 5564 4196 5572 4204
rect 5628 4156 5636 4164
rect 5596 4096 5604 4104
rect 5580 3936 5588 3944
rect 5564 3896 5572 3904
rect 5356 3836 5364 3844
rect 5276 3776 5284 3784
rect 5308 3776 5316 3784
rect 5372 3776 5380 3784
rect 5052 3736 5060 3744
rect 5084 3736 5092 3744
rect 5116 3736 5124 3744
rect 5196 3736 5204 3744
rect 5260 3736 5268 3744
rect 5020 3676 5028 3684
rect 5228 3716 5236 3724
rect 5164 3656 5172 3664
rect 5180 3656 5188 3664
rect 5084 3636 5092 3644
rect 5116 3596 5124 3604
rect 5196 3576 5204 3584
rect 5196 3536 5204 3544
rect 5228 3536 5236 3544
rect 5212 3516 5220 3524
rect 5036 3496 5044 3504
rect 5084 3496 5092 3504
rect 5004 3436 5012 3444
rect 5068 3416 5076 3424
rect 5116 3416 5124 3424
rect 5004 3376 5012 3384
rect 5052 3376 5060 3384
rect 4924 3356 4932 3364
rect 5068 3356 5076 3364
rect 5100 3356 5108 3364
rect 4892 3336 4900 3344
rect 4940 3336 4948 3344
rect 4972 3336 4980 3344
rect 5020 3336 5028 3344
rect 5052 3336 5060 3344
rect 5068 3336 5076 3344
rect 4892 3296 4900 3304
rect 4972 3276 4980 3284
rect 4924 3256 4932 3264
rect 5020 3256 5028 3264
rect 4988 3136 4996 3144
rect 4876 3056 4884 3064
rect 4860 3016 4868 3024
rect 5004 3056 5012 3064
rect 4940 3036 4948 3044
rect 4924 2996 4932 3004
rect 4956 2976 4964 2984
rect 4764 2896 4772 2904
rect 4812 2896 4820 2904
rect 4828 2896 4836 2904
rect 4540 2876 4548 2884
rect 4716 2876 4724 2884
rect 4524 2796 4532 2804
rect 4508 2776 4516 2784
rect 4412 2736 4420 2744
rect 4428 2736 4436 2744
rect 4364 2716 4372 2724
rect 4428 2716 4436 2724
rect 4460 2716 4468 2724
rect 4348 2696 4356 2704
rect 4524 2716 4532 2724
rect 4412 2696 4420 2704
rect 4492 2696 4500 2704
rect 4172 2676 4180 2684
rect 4396 2676 4404 2684
rect 4396 2656 4404 2664
rect 4140 2636 4148 2644
rect 4156 2636 4164 2644
rect 4204 2636 4212 2644
rect 4428 2636 4436 2644
rect 4140 2616 4148 2624
rect 4124 2496 4132 2504
rect 4124 2436 4132 2444
rect 3756 2176 3764 2184
rect 3852 2176 3860 2184
rect 3916 2176 3924 2184
rect 3996 2176 4004 2184
rect 4108 2176 4116 2184
rect 3740 2156 3748 2164
rect 3708 2136 3716 2144
rect 3740 2096 3748 2104
rect 3740 2056 3748 2064
rect 3708 2036 3716 2044
rect 3724 2016 3732 2024
rect 3708 1916 3716 1924
rect 3740 1916 3748 1924
rect 3708 1896 3716 1904
rect 3740 1896 3748 1904
rect 3724 1856 3732 1864
rect 3692 1776 3700 1784
rect 3676 1756 3684 1764
rect 3708 1756 3716 1764
rect 3692 1736 3700 1744
rect 3676 1696 3684 1704
rect 3676 1556 3684 1564
rect 3724 1536 3732 1544
rect 3660 1476 3668 1484
rect 3644 1436 3652 1444
rect 3644 1416 3652 1424
rect 3628 1376 3636 1384
rect 3628 1356 3636 1364
rect 3596 1336 3604 1344
rect 3580 1196 3588 1204
rect 3596 1196 3604 1204
rect 3820 2156 3828 2164
rect 3900 2156 3908 2164
rect 3772 2116 3780 2124
rect 3772 2096 3780 2104
rect 3980 2156 3988 2164
rect 3948 2136 3956 2144
rect 3884 2116 3892 2124
rect 3868 2076 3876 2084
rect 3900 2076 3908 2084
rect 3788 2036 3796 2044
rect 3820 1936 3828 1944
rect 3868 1916 3876 1924
rect 3788 1876 3796 1884
rect 3836 1876 3844 1884
rect 3820 1776 3828 1784
rect 3852 1776 3860 1784
rect 3868 1776 3876 1784
rect 3916 2036 3924 2044
rect 4012 2156 4020 2164
rect 4028 2136 4036 2144
rect 4012 2116 4020 2124
rect 4076 2116 4084 2124
rect 4108 2116 4116 2124
rect 4108 2076 4116 2084
rect 4092 2036 4100 2044
rect 4140 2316 4148 2324
rect 4124 1996 4132 2004
rect 4140 1996 4148 2004
rect 4108 1976 4116 1984
rect 4044 1956 4052 1964
rect 4060 1956 4068 1964
rect 3932 1876 3940 1884
rect 3996 1876 4004 1884
rect 3948 1856 3956 1864
rect 3980 1856 3988 1864
rect 4188 2596 4196 2604
rect 4220 2596 4228 2604
rect 4588 2856 4596 2864
rect 4638 2806 4646 2814
rect 4652 2806 4660 2814
rect 4666 2806 4674 2814
rect 4764 2796 4772 2804
rect 4556 2696 4564 2704
rect 4604 2696 4612 2704
rect 4572 2676 4580 2684
rect 4652 2676 4660 2684
rect 4572 2636 4580 2644
rect 4684 2596 4692 2604
rect 4444 2576 4452 2584
rect 4508 2576 4516 2584
rect 4268 2556 4276 2564
rect 4380 2556 4388 2564
rect 4396 2556 4404 2564
rect 4252 2536 4260 2544
rect 4412 2536 4420 2544
rect 4300 2516 4308 2524
rect 4252 2496 4260 2504
rect 4284 2496 4292 2504
rect 4332 2496 4340 2504
rect 4428 2496 4436 2504
rect 4236 2476 4244 2484
rect 4316 2476 4324 2484
rect 4396 2476 4404 2484
rect 4268 2456 4276 2464
rect 4284 2456 4292 2464
rect 4380 2456 4388 2464
rect 4220 2396 4228 2404
rect 4252 2396 4260 2404
rect 4172 2376 4180 2384
rect 4204 2376 4212 2384
rect 4188 2316 4196 2324
rect 4316 2416 4324 2424
rect 4268 2296 4276 2304
rect 4364 2376 4372 2384
rect 4380 2376 4388 2384
rect 4348 2316 4356 2324
rect 4332 2296 4340 2304
rect 4412 2456 4420 2464
rect 4652 2556 4660 2564
rect 4476 2536 4484 2544
rect 4524 2536 4532 2544
rect 4556 2536 4564 2544
rect 4588 2536 4596 2544
rect 4604 2536 4612 2544
rect 4460 2516 4468 2524
rect 4572 2496 4580 2504
rect 4572 2436 4580 2444
rect 4556 2396 4564 2404
rect 4796 2716 4804 2724
rect 4796 2696 4804 2704
rect 4748 2676 4756 2684
rect 5100 3236 5108 3244
rect 5084 3216 5092 3224
rect 5068 3196 5076 3204
rect 5036 3096 5044 3104
rect 5068 3056 5076 3064
rect 5116 3196 5124 3204
rect 5116 3176 5124 3184
rect 5100 2976 5108 2984
rect 5036 2916 5044 2924
rect 5084 2916 5092 2924
rect 5004 2876 5012 2884
rect 4988 2836 4996 2844
rect 5020 2836 5028 2844
rect 4860 2776 4868 2784
rect 4892 2756 4900 2764
rect 4908 2756 4916 2764
rect 4828 2696 4836 2704
rect 4844 2696 4852 2704
rect 4812 2676 4820 2684
rect 4876 2636 4884 2644
rect 4716 2596 4724 2604
rect 4700 2556 4708 2564
rect 4684 2496 4692 2504
rect 4636 2476 4644 2484
rect 4604 2416 4612 2424
rect 4638 2406 4646 2414
rect 4652 2406 4660 2414
rect 4666 2406 4674 2414
rect 4700 2396 4708 2404
rect 4444 2376 4452 2384
rect 4588 2376 4596 2384
rect 4652 2376 4660 2384
rect 4748 2436 4756 2444
rect 4604 2336 4612 2344
rect 4428 2316 4436 2324
rect 4492 2316 4500 2324
rect 4636 2316 4644 2324
rect 4508 2296 4516 2304
rect 4668 2296 4676 2304
rect 4428 2276 4436 2284
rect 4572 2276 4580 2284
rect 4220 2256 4228 2264
rect 4316 2256 4324 2264
rect 4540 2256 4548 2264
rect 4588 2256 4596 2264
rect 4220 2196 4228 2204
rect 4236 2196 4244 2204
rect 4188 2176 4196 2184
rect 4220 2176 4228 2184
rect 4236 2176 4244 2184
rect 4172 2136 4180 2144
rect 4460 2236 4468 2244
rect 4268 2216 4276 2224
rect 4444 2196 4452 2204
rect 4508 2196 4516 2204
rect 4412 2176 4420 2184
rect 4476 2176 4484 2184
rect 4268 2136 4276 2144
rect 4300 2136 4308 2144
rect 4348 2136 4356 2144
rect 4396 2136 4404 2144
rect 4204 2116 4212 2124
rect 4252 2116 4260 2124
rect 4188 2056 4196 2064
rect 4460 2136 4468 2144
rect 4508 2136 4516 2144
rect 4604 2136 4612 2144
rect 4396 2116 4404 2124
rect 4444 2116 4452 2124
rect 4284 2036 4292 2044
rect 4716 2376 4724 2384
rect 4700 2276 4708 2284
rect 4764 2416 4772 2424
rect 4844 2576 4852 2584
rect 4812 2536 4820 2544
rect 4828 2536 4836 2544
rect 4780 2376 4788 2384
rect 4924 2676 4932 2684
rect 5068 2876 5076 2884
rect 5052 2796 5060 2804
rect 4972 2776 4980 2784
rect 5004 2776 5012 2784
rect 5100 2776 5108 2784
rect 5004 2756 5012 2764
rect 5068 2756 5076 2764
rect 5100 2756 5108 2764
rect 4956 2716 4964 2724
rect 4972 2716 4980 2724
rect 5020 2696 5028 2704
rect 4988 2676 4996 2684
rect 4940 2636 4948 2644
rect 4956 2636 4964 2644
rect 5084 2716 5092 2724
rect 5068 2696 5076 2704
rect 5052 2676 5060 2684
rect 5036 2636 5044 2644
rect 4940 2536 4948 2544
rect 5004 2536 5012 2544
rect 5036 2536 5044 2544
rect 4828 2476 4836 2484
rect 4860 2476 4868 2484
rect 4812 2416 4820 2424
rect 4828 2416 4836 2424
rect 4924 2476 4932 2484
rect 4972 2476 4980 2484
rect 4828 2376 4836 2384
rect 4876 2376 4884 2384
rect 4940 2376 4948 2384
rect 4956 2376 4964 2384
rect 4764 2316 4772 2324
rect 4748 2296 4756 2304
rect 4780 2296 4788 2304
rect 4764 2276 4772 2284
rect 4732 2236 4740 2244
rect 4748 2236 4756 2244
rect 4716 2216 4724 2224
rect 4764 2216 4772 2224
rect 4956 2316 4964 2324
rect 4812 2276 4820 2284
rect 4844 2276 4852 2284
rect 4796 2236 4804 2244
rect 4716 2156 4724 2164
rect 4732 2156 4740 2164
rect 4524 2116 4532 2124
rect 4572 2116 4580 2124
rect 4348 2076 4356 2084
rect 4508 2076 4516 2084
rect 4540 2076 4548 2084
rect 4540 2056 4548 2064
rect 4556 2056 4564 2064
rect 4316 2036 4324 2044
rect 4380 2036 4388 2044
rect 4396 2036 4404 2044
rect 4300 1996 4308 2004
rect 4348 2016 4356 2024
rect 4284 1916 4292 1924
rect 4332 1916 4340 1924
rect 4348 1916 4356 1924
rect 4380 1916 4388 1924
rect 4172 1896 4180 1904
rect 4028 1876 4036 1884
rect 4076 1876 4084 1884
rect 4108 1876 4116 1884
rect 4124 1876 4132 1884
rect 4156 1856 4164 1864
rect 3916 1816 3924 1824
rect 3964 1816 3972 1824
rect 4012 1816 4020 1824
rect 4060 1816 4068 1824
rect 4140 1796 4148 1804
rect 4156 1796 4164 1804
rect 4060 1776 4068 1784
rect 4140 1776 4148 1784
rect 3900 1736 3908 1744
rect 3788 1656 3796 1664
rect 3772 1596 3780 1604
rect 3756 1556 3764 1564
rect 3868 1676 3876 1684
rect 3948 1736 3956 1744
rect 4012 1736 4020 1744
rect 3852 1636 3860 1644
rect 3932 1636 3940 1644
rect 3884 1616 3892 1624
rect 4092 1676 4100 1684
rect 4028 1656 4036 1664
rect 4124 1736 4132 1744
rect 4124 1676 4132 1684
rect 4204 1896 4212 1904
rect 4204 1876 4212 1884
rect 4252 1876 4260 1884
rect 4220 1856 4228 1864
rect 4332 1856 4340 1864
rect 4412 1956 4420 1964
rect 4428 1916 4436 1924
rect 4444 1896 4452 1904
rect 4188 1836 4196 1844
rect 4284 1836 4292 1844
rect 4364 1836 4372 1844
rect 4220 1816 4228 1824
rect 4188 1796 4196 1804
rect 3996 1636 4004 1644
rect 4108 1636 4116 1644
rect 3964 1616 3972 1624
rect 4124 1616 4132 1624
rect 3804 1596 3812 1604
rect 3932 1596 3940 1604
rect 3948 1596 3956 1604
rect 3804 1576 3812 1584
rect 3916 1576 3924 1584
rect 3852 1556 3860 1564
rect 3868 1556 3876 1564
rect 3804 1536 3812 1544
rect 3772 1516 3780 1524
rect 3900 1516 3908 1524
rect 3980 1596 3988 1604
rect 4076 1596 4084 1604
rect 3948 1516 3956 1524
rect 4060 1556 4068 1564
rect 4028 1516 4036 1524
rect 4044 1516 4052 1524
rect 3980 1476 3988 1484
rect 3804 1436 3812 1444
rect 3868 1436 3876 1444
rect 3740 1396 3748 1404
rect 3772 1376 3780 1384
rect 3708 1356 3716 1364
rect 3916 1416 3924 1424
rect 3932 1416 3940 1424
rect 3788 1356 3796 1364
rect 3916 1356 3924 1364
rect 3676 1316 3684 1324
rect 3692 1316 3700 1324
rect 3724 1316 3732 1324
rect 3756 1316 3764 1324
rect 3644 1276 3652 1284
rect 3660 1276 3668 1284
rect 3708 1276 3716 1284
rect 3660 1236 3668 1244
rect 3644 1196 3652 1204
rect 3564 1176 3572 1184
rect 3564 1156 3572 1164
rect 3612 1156 3620 1164
rect 3628 1156 3636 1164
rect 3548 1136 3556 1144
rect 3532 1116 3540 1124
rect 3180 1076 3188 1084
rect 3212 1076 3220 1084
rect 3260 1076 3268 1084
rect 3292 1076 3300 1084
rect 3324 1076 3332 1084
rect 3356 1076 3364 1084
rect 3324 1056 3332 1064
rect 3068 1036 3076 1044
rect 3180 1016 3188 1024
rect 3118 1006 3126 1014
rect 3132 1006 3140 1014
rect 3146 1006 3154 1014
rect 3084 996 3092 1004
rect 3260 996 3268 1004
rect 3276 996 3284 1004
rect 3116 956 3124 964
rect 3228 916 3236 924
rect 3276 916 3284 924
rect 3292 916 3300 924
rect 2940 876 2948 884
rect 3036 876 3044 884
rect 3052 876 3060 884
rect 3260 876 3268 884
rect 2924 856 2932 864
rect 2764 736 2772 744
rect 2844 736 2852 744
rect 2780 716 2788 724
rect 2796 696 2804 704
rect 2876 696 2884 704
rect 2956 816 2964 824
rect 3084 816 3092 824
rect 3036 756 3044 764
rect 2924 696 2932 704
rect 2956 696 2964 704
rect 3052 696 3060 704
rect 2812 676 2820 684
rect 2844 676 2852 684
rect 2908 676 2916 684
rect 2972 676 2980 684
rect 3020 676 3028 684
rect 2828 656 2836 664
rect 2972 656 2980 664
rect 3068 656 3076 664
rect 2812 636 2820 644
rect 2796 596 2804 604
rect 2732 576 2740 584
rect 2764 576 2772 584
rect 2604 556 2612 564
rect 2572 536 2580 544
rect 2604 536 2612 544
rect 2780 536 2788 544
rect 2556 516 2564 524
rect 2524 496 2532 504
rect 2716 476 2724 484
rect 2764 476 2772 484
rect 2620 456 2628 464
rect 2732 456 2740 464
rect 2892 596 2900 604
rect 2844 556 2852 564
rect 2860 536 2868 544
rect 2876 536 2884 544
rect 2940 536 2948 544
rect 3004 536 3012 544
rect 3036 536 3044 544
rect 3020 516 3028 524
rect 3068 516 3076 524
rect 2956 476 2964 484
rect 2892 456 2900 464
rect 2812 436 2820 444
rect 2540 416 2548 424
rect 2940 436 2948 444
rect 3004 396 3012 404
rect 2444 376 2452 384
rect 2588 356 2596 364
rect 2796 336 2804 344
rect 2844 336 2852 344
rect 2908 336 2916 344
rect 2428 316 2436 324
rect 2476 316 2484 324
rect 2492 316 2500 324
rect 2636 316 2644 324
rect 2716 316 2724 324
rect 2764 316 2772 324
rect 2460 296 2468 304
rect 2364 276 2372 284
rect 2428 276 2436 284
rect 2444 236 2452 244
rect 2412 216 2420 224
rect 2332 156 2340 164
rect 2380 156 2388 164
rect 2188 136 2196 144
rect 2188 116 2196 124
rect 2156 16 2164 24
rect 2236 116 2244 124
rect 2348 116 2356 124
rect 2332 16 2340 24
rect 2556 296 2564 304
rect 2604 276 2612 284
rect 2652 296 2660 304
rect 2812 316 2820 324
rect 2812 296 2820 304
rect 2652 276 2660 284
rect 2860 316 2868 324
rect 2892 296 2900 304
rect 3068 316 3076 324
rect 2924 276 2932 284
rect 2636 256 2644 264
rect 2748 256 2756 264
rect 2764 236 2772 244
rect 2828 216 2836 224
rect 2764 196 2772 204
rect 2988 236 2996 244
rect 3036 236 3044 244
rect 3164 696 3172 704
rect 3212 796 3220 804
rect 3196 736 3204 744
rect 3308 776 3316 784
rect 3340 776 3348 784
rect 3260 676 3268 684
rect 3260 656 3268 664
rect 3372 1056 3380 1064
rect 3388 1056 3396 1064
rect 3420 1036 3428 1044
rect 3436 1036 3444 1044
rect 3580 1136 3588 1144
rect 3596 1116 3604 1124
rect 3884 1316 3892 1324
rect 3820 1276 3828 1284
rect 3852 1276 3860 1284
rect 3788 1236 3796 1244
rect 3868 1216 3876 1224
rect 3740 1196 3748 1204
rect 3756 1196 3764 1204
rect 3756 1176 3764 1184
rect 3756 1156 3764 1164
rect 3692 1136 3700 1144
rect 3740 1136 3748 1144
rect 3660 1116 3668 1124
rect 3724 1116 3732 1124
rect 3772 1116 3780 1124
rect 3644 1096 3652 1104
rect 3708 1096 3716 1104
rect 3500 1036 3508 1044
rect 3548 1036 3556 1044
rect 3468 1016 3476 1024
rect 3484 1016 3492 1024
rect 3452 996 3460 1004
rect 3388 976 3396 984
rect 3372 956 3380 964
rect 3436 956 3444 964
rect 3452 936 3460 944
rect 3564 1016 3572 1024
rect 3580 1016 3588 1024
rect 3564 936 3572 944
rect 3836 1096 3844 1104
rect 3772 976 3780 984
rect 3692 956 3700 964
rect 3836 1016 3844 1024
rect 3852 1016 3860 1024
rect 3900 1276 3908 1284
rect 3900 1236 3908 1244
rect 3916 1216 3924 1224
rect 3900 1176 3908 1184
rect 3916 1176 3924 1184
rect 3900 1096 3908 1104
rect 3980 1376 3988 1384
rect 3964 1356 3972 1364
rect 4028 1476 4036 1484
rect 4092 1556 4100 1564
rect 4108 1556 4116 1564
rect 4172 1556 4180 1564
rect 4124 1536 4132 1544
rect 4108 1496 4116 1504
rect 4364 1796 4372 1804
rect 4316 1776 4324 1784
rect 4300 1716 4308 1724
rect 4204 1656 4212 1664
rect 4220 1556 4228 1564
rect 4300 1696 4308 1704
rect 4332 1696 4340 1704
rect 4268 1676 4276 1684
rect 4252 1576 4260 1584
rect 4236 1516 4244 1524
rect 4268 1556 4276 1564
rect 4284 1496 4292 1504
rect 4140 1476 4148 1484
rect 4188 1476 4196 1484
rect 4252 1476 4260 1484
rect 4284 1456 4292 1464
rect 4156 1396 4164 1404
rect 4060 1356 4068 1364
rect 4108 1356 4116 1364
rect 4140 1356 4148 1364
rect 3948 1316 3956 1324
rect 3996 1316 4004 1324
rect 4028 1296 4036 1304
rect 4028 1196 4036 1204
rect 4012 1176 4020 1184
rect 3996 1156 4004 1164
rect 4108 1336 4116 1344
rect 4172 1336 4180 1344
rect 4156 1316 4164 1324
rect 4284 1416 4292 1424
rect 4204 1396 4212 1404
rect 4252 1356 4260 1364
rect 4220 1336 4228 1344
rect 4204 1316 4212 1324
rect 4252 1296 4260 1304
rect 4284 1336 4292 1344
rect 4188 1276 4196 1284
rect 4076 1136 4084 1144
rect 4348 1676 4356 1684
rect 4364 1576 4372 1584
rect 4332 1516 4340 1524
rect 4316 1476 4324 1484
rect 4348 1416 4356 1424
rect 4316 1376 4324 1384
rect 4332 1376 4340 1384
rect 4332 1316 4340 1324
rect 4316 1276 4324 1284
rect 4252 1256 4260 1264
rect 4300 1256 4308 1264
rect 4172 1216 4180 1224
rect 4204 1216 4212 1224
rect 4204 1196 4212 1204
rect 4364 1236 4372 1244
rect 4428 1876 4436 1884
rect 4460 1876 4468 1884
rect 4492 1896 4500 1904
rect 4540 1876 4548 1884
rect 4556 1876 4564 1884
rect 4476 1856 4484 1864
rect 4508 1856 4516 1864
rect 4396 1796 4404 1804
rect 4460 1776 4468 1784
rect 4428 1756 4436 1764
rect 4476 1756 4484 1764
rect 4396 1736 4404 1744
rect 4412 1676 4420 1684
rect 4396 1656 4404 1664
rect 4396 1556 4404 1564
rect 4588 2076 4596 2084
rect 4604 2076 4612 2084
rect 4620 2056 4628 2064
rect 4638 2006 4646 2014
rect 4652 2006 4660 2014
rect 4666 2006 4674 2014
rect 4732 2136 4740 2144
rect 4716 2036 4724 2044
rect 4828 2256 4836 2264
rect 4956 2256 4964 2264
rect 4940 2236 4948 2244
rect 4892 2216 4900 2224
rect 4844 2156 4852 2164
rect 4812 2116 4820 2124
rect 4604 1956 4612 1964
rect 4620 1916 4628 1924
rect 4588 1836 4596 1844
rect 4652 1836 4660 1844
rect 4572 1796 4580 1804
rect 4524 1736 4532 1744
rect 4524 1716 4532 1724
rect 4428 1636 4436 1644
rect 4428 1576 4436 1584
rect 4412 1516 4420 1524
rect 4412 1436 4420 1444
rect 4380 1216 4388 1224
rect 4364 1176 4372 1184
rect 4588 1736 4596 1744
rect 4684 1716 4692 1724
rect 4700 1716 4708 1724
rect 4764 2016 4772 2024
rect 4828 1996 4836 2004
rect 4860 2096 4868 2104
rect 4844 1956 4852 1964
rect 4828 1916 4836 1924
rect 4812 1896 4820 1904
rect 4732 1876 4740 1884
rect 4780 1856 4788 1864
rect 4748 1836 4756 1844
rect 4764 1776 4772 1784
rect 4572 1696 4580 1704
rect 4716 1696 4724 1704
rect 4732 1696 4740 1704
rect 4540 1656 4548 1664
rect 4476 1596 4484 1604
rect 4460 1556 4468 1564
rect 4460 1536 4468 1544
rect 4444 1476 4452 1484
rect 4444 1356 4452 1364
rect 4428 1316 4436 1324
rect 4460 1276 4468 1284
rect 4492 1516 4500 1524
rect 4508 1516 4516 1524
rect 4638 1606 4646 1614
rect 4652 1606 4660 1614
rect 4666 1606 4674 1614
rect 4556 1576 4564 1584
rect 4652 1576 4660 1584
rect 4572 1516 4580 1524
rect 4588 1516 4596 1524
rect 4524 1456 4532 1464
rect 4876 1956 4884 1964
rect 4956 2216 4964 2224
rect 5020 2396 5028 2404
rect 4988 2376 4996 2384
rect 5052 2456 5060 2464
rect 5036 2336 5044 2344
rect 5244 3496 5252 3504
rect 5340 3616 5348 3624
rect 5548 3856 5556 3864
rect 5500 3816 5508 3824
rect 5516 3776 5524 3784
rect 5420 3736 5428 3744
rect 5452 3736 5460 3744
rect 5468 3740 5476 3744
rect 5468 3736 5476 3740
rect 5404 3716 5412 3724
rect 5436 3676 5444 3684
rect 5452 3676 5460 3684
rect 5388 3636 5396 3644
rect 5420 3636 5428 3644
rect 5356 3596 5364 3604
rect 5276 3536 5284 3544
rect 5404 3516 5412 3524
rect 5308 3496 5316 3504
rect 5324 3496 5332 3504
rect 5196 3476 5204 3484
rect 5260 3476 5268 3484
rect 5212 3456 5220 3464
rect 5244 3456 5252 3464
rect 5164 3416 5172 3424
rect 5292 3456 5300 3464
rect 5132 3096 5140 3104
rect 5132 2996 5140 3004
rect 5228 3316 5236 3324
rect 5212 3276 5220 3284
rect 5180 3236 5188 3244
rect 5164 3116 5172 3124
rect 5292 3296 5300 3304
rect 5260 3236 5268 3244
rect 5228 3096 5236 3104
rect 5164 3076 5172 3084
rect 5212 3056 5220 3064
rect 5180 3036 5188 3044
rect 5292 3156 5300 3164
rect 5244 3076 5252 3084
rect 5292 3056 5300 3064
rect 5324 3436 5332 3444
rect 5372 3436 5380 3444
rect 5404 3416 5412 3424
rect 5356 3356 5364 3364
rect 5324 3296 5332 3304
rect 5340 3296 5348 3304
rect 5484 3636 5492 3644
rect 5548 3756 5556 3764
rect 5532 3636 5540 3644
rect 5484 3616 5492 3624
rect 5516 3616 5524 3624
rect 5452 3536 5460 3544
rect 5436 3496 5444 3504
rect 5468 3516 5476 3524
rect 5436 3456 5444 3464
rect 5452 3336 5460 3344
rect 5436 3316 5444 3324
rect 5420 3216 5428 3224
rect 5372 3136 5380 3144
rect 5324 3116 5332 3124
rect 5452 3296 5460 3304
rect 5468 3096 5476 3104
rect 5340 3076 5348 3084
rect 5404 3016 5412 3024
rect 5308 2996 5316 3004
rect 5212 2956 5220 2964
rect 5228 2956 5236 2964
rect 5164 2916 5172 2924
rect 5196 2816 5204 2824
rect 5212 2816 5220 2824
rect 5148 2776 5156 2784
rect 5180 2776 5188 2784
rect 5196 2776 5204 2784
rect 5132 2756 5140 2764
rect 5164 2716 5172 2724
rect 5196 2756 5204 2764
rect 5212 2756 5220 2764
rect 5116 2636 5124 2644
rect 5180 2636 5188 2644
rect 5148 2616 5156 2624
rect 5164 2596 5172 2604
rect 5148 2556 5156 2564
rect 5132 2536 5140 2544
rect 5116 2496 5124 2504
rect 5100 2476 5108 2484
rect 5116 2456 5124 2464
rect 5116 2396 5124 2404
rect 5084 2316 5092 2324
rect 5100 2316 5108 2324
rect 5004 2276 5012 2284
rect 4988 2256 4996 2264
rect 5020 2256 5028 2264
rect 4940 2156 4948 2164
rect 4988 2176 4996 2184
rect 5020 2176 5028 2184
rect 4972 2156 4980 2164
rect 5052 2276 5060 2284
rect 5084 2256 5092 2264
rect 5212 2616 5220 2624
rect 5372 2976 5380 2984
rect 5356 2916 5364 2924
rect 5452 2976 5460 2984
rect 5388 2896 5396 2904
rect 5292 2836 5300 2844
rect 5356 2836 5364 2844
rect 5276 2776 5284 2784
rect 5244 2756 5252 2764
rect 5420 2876 5428 2884
rect 5388 2816 5396 2824
rect 5404 2816 5412 2824
rect 5244 2716 5252 2724
rect 5276 2736 5284 2744
rect 5292 2736 5300 2744
rect 5436 2656 5444 2664
rect 5308 2636 5316 2644
rect 5292 2596 5300 2604
rect 5404 2596 5412 2604
rect 5260 2576 5268 2584
rect 5212 2556 5220 2564
rect 5228 2556 5236 2564
rect 5308 2556 5316 2564
rect 5372 2556 5380 2564
rect 5244 2536 5252 2544
rect 5276 2536 5284 2544
rect 5244 2476 5252 2484
rect 5276 2476 5284 2484
rect 5276 2376 5284 2384
rect 5180 2336 5188 2344
rect 5276 2336 5284 2344
rect 5164 2316 5172 2324
rect 5212 2316 5220 2324
rect 5132 2296 5140 2304
rect 5324 2536 5332 2544
rect 5388 2516 5396 2524
rect 5436 2556 5444 2564
rect 5420 2536 5428 2544
rect 5436 2516 5444 2524
rect 5340 2476 5348 2484
rect 5468 2856 5476 2864
rect 5516 3556 5524 3564
rect 5500 3496 5508 3504
rect 5532 3496 5540 3504
rect 5644 4116 5652 4124
rect 5852 4596 5860 4604
rect 5836 4556 5844 4564
rect 5932 4896 5940 4904
rect 5916 4876 5924 4884
rect 6140 5756 6148 5764
rect 6172 5756 6180 5764
rect 6124 5696 6132 5704
rect 6172 5696 6180 5704
rect 6188 5676 6196 5684
rect 6156 5496 6164 5504
rect 6172 5476 6180 5484
rect 6108 5376 6116 5384
rect 6172 5376 6180 5384
rect 6236 5536 6244 5544
rect 6220 5356 6228 5364
rect 6220 5336 6228 5344
rect 6188 5316 6196 5324
rect 6188 5216 6196 5224
rect 6252 5236 6260 5244
rect 6252 5216 6260 5224
rect 6204 5136 6212 5144
rect 6188 5076 6196 5084
rect 6060 5056 6068 5064
rect 6220 5096 6228 5104
rect 6076 5036 6084 5044
rect 5980 4976 5988 4984
rect 5996 4976 6004 4984
rect 5964 4956 5972 4964
rect 5964 4896 5972 4904
rect 5948 4856 5956 4864
rect 5900 4776 5908 4784
rect 5884 4676 5892 4684
rect 5932 4776 5940 4784
rect 5932 4756 5940 4764
rect 5948 4716 5956 4724
rect 5884 4636 5892 4644
rect 5900 4596 5908 4604
rect 6028 4956 6036 4964
rect 6108 4996 6116 5004
rect 6172 4936 6180 4944
rect 6220 5056 6228 5064
rect 6236 5016 6244 5024
rect 5996 4856 6004 4864
rect 5980 4796 5988 4804
rect 5980 4696 5988 4704
rect 6044 4836 6052 4844
rect 6060 4836 6068 4844
rect 6140 4836 6148 4844
rect 6060 4796 6068 4804
rect 6060 4756 6068 4764
rect 6044 4716 6052 4724
rect 6156 4736 6164 4744
rect 6076 4716 6084 4724
rect 6108 4716 6116 4724
rect 6028 4676 6036 4684
rect 6012 4656 6020 4664
rect 6028 4656 6036 4664
rect 5964 4616 5972 4624
rect 5980 4576 5988 4584
rect 5836 4536 5844 4544
rect 5868 4536 5876 4544
rect 5740 4476 5748 4484
rect 5788 4476 5796 4484
rect 5820 4336 5828 4344
rect 5868 4516 5876 4524
rect 5964 4536 5972 4544
rect 5996 4540 6004 4544
rect 5996 4536 6004 4540
rect 5916 4516 5924 4524
rect 5852 4476 5860 4484
rect 5724 4296 5732 4304
rect 5740 4296 5748 4304
rect 5804 4296 5812 4304
rect 5836 4296 5844 4304
rect 5900 4496 5908 4504
rect 5932 4476 5940 4484
rect 5916 4356 5924 4364
rect 5868 4296 5876 4304
rect 5916 4296 5924 4304
rect 5836 4276 5844 4284
rect 5852 4276 5860 4284
rect 5740 4256 5748 4264
rect 5708 4216 5716 4224
rect 5740 4216 5748 4224
rect 5676 4156 5684 4164
rect 5692 4156 5700 4164
rect 5724 4156 5732 4164
rect 5628 4096 5636 4104
rect 5660 4096 5668 4104
rect 5660 4076 5668 4084
rect 5708 4136 5716 4144
rect 5692 4076 5700 4084
rect 5676 4056 5684 4064
rect 5676 4036 5684 4044
rect 5756 4156 5764 4164
rect 5756 4116 5764 4124
rect 5724 4056 5732 4064
rect 5660 3916 5668 3924
rect 5660 3896 5668 3904
rect 5644 3876 5652 3884
rect 5612 3856 5620 3864
rect 5596 3776 5604 3784
rect 5612 3756 5620 3764
rect 5660 3796 5668 3804
rect 5740 3936 5748 3944
rect 5708 3916 5716 3924
rect 5708 3876 5716 3884
rect 5724 3876 5732 3884
rect 5692 3856 5700 3864
rect 5724 3816 5732 3824
rect 5692 3796 5700 3804
rect 5660 3776 5668 3784
rect 5596 3736 5604 3744
rect 5612 3736 5620 3744
rect 5628 3736 5636 3744
rect 5580 3716 5588 3724
rect 5564 3476 5572 3484
rect 5532 3456 5540 3464
rect 5532 3436 5540 3444
rect 5644 3696 5652 3704
rect 5708 3756 5716 3764
rect 5708 3736 5716 3744
rect 5628 3656 5636 3664
rect 5612 3596 5620 3604
rect 5596 3516 5604 3524
rect 5580 3396 5588 3404
rect 5548 3356 5556 3364
rect 5676 3656 5684 3664
rect 5660 3556 5668 3564
rect 5628 3396 5636 3404
rect 5644 3376 5652 3384
rect 5628 3356 5636 3364
rect 5660 3356 5668 3364
rect 5516 3336 5524 3344
rect 5612 3336 5620 3344
rect 5500 3316 5508 3324
rect 5580 3316 5588 3324
rect 5580 3296 5588 3304
rect 5516 3196 5524 3204
rect 5548 3196 5556 3204
rect 5500 3116 5508 3124
rect 5532 3116 5540 3124
rect 5500 3076 5508 3084
rect 5516 3036 5524 3044
rect 5564 3056 5572 3064
rect 5532 2956 5540 2964
rect 5548 2956 5556 2964
rect 5612 3156 5620 3164
rect 5644 3336 5652 3344
rect 5644 3316 5652 3324
rect 5724 3576 5732 3584
rect 5836 4256 5844 4264
rect 5788 4216 5796 4224
rect 5852 4236 5860 4244
rect 5820 4176 5828 4184
rect 5804 4136 5812 4144
rect 5836 4136 5844 4144
rect 5884 4276 5892 4284
rect 5932 4276 5940 4284
rect 5932 4256 5940 4264
rect 5900 4216 5908 4224
rect 5788 4096 5796 4104
rect 5836 4096 5844 4104
rect 5772 3996 5780 4004
rect 5772 3796 5780 3804
rect 5772 3756 5780 3764
rect 5756 3736 5764 3744
rect 5820 3996 5828 4004
rect 5804 3976 5812 3984
rect 5836 3936 5844 3944
rect 5820 3896 5828 3904
rect 5884 4076 5892 4084
rect 5868 4056 5876 4064
rect 5868 4036 5876 4044
rect 5916 4036 5924 4044
rect 5900 4016 5908 4024
rect 5884 3996 5892 4004
rect 5900 3996 5908 4004
rect 5868 3976 5876 3984
rect 5884 3936 5892 3944
rect 5948 4236 5956 4244
rect 5980 4476 5988 4484
rect 5980 4356 5988 4364
rect 6012 4356 6020 4364
rect 5948 4076 5956 4084
rect 5964 4056 5972 4064
rect 5932 3996 5940 4004
rect 5948 3996 5956 4004
rect 5916 3956 5924 3964
rect 5884 3896 5892 3904
rect 5820 3816 5828 3824
rect 5820 3796 5828 3804
rect 5804 3756 5812 3764
rect 5820 3736 5828 3744
rect 5756 3716 5764 3724
rect 5788 3716 5796 3724
rect 5804 3696 5812 3704
rect 5788 3676 5796 3684
rect 5772 3596 5780 3604
rect 5788 3596 5796 3604
rect 5788 3576 5796 3584
rect 5740 3556 5748 3564
rect 5756 3536 5764 3544
rect 5692 3516 5700 3524
rect 5740 3516 5748 3524
rect 5692 3456 5700 3464
rect 5788 3516 5796 3524
rect 5772 3476 5780 3484
rect 5740 3416 5748 3424
rect 5756 3396 5764 3404
rect 5788 3456 5796 3464
rect 5788 3416 5796 3424
rect 5708 3336 5716 3344
rect 5740 3340 5748 3344
rect 5740 3336 5748 3340
rect 5676 3256 5684 3264
rect 5660 3196 5668 3204
rect 5756 3276 5764 3284
rect 5788 3256 5796 3264
rect 5740 3236 5748 3244
rect 5708 3156 5716 3164
rect 5644 3136 5652 3144
rect 5628 3096 5636 3104
rect 5612 3076 5620 3084
rect 5580 3016 5588 3024
rect 5596 3016 5604 3024
rect 5564 2936 5572 2944
rect 5564 2896 5572 2904
rect 5660 3116 5668 3124
rect 5676 3116 5684 3124
rect 5660 3096 5668 3104
rect 5628 2976 5636 2984
rect 5692 3056 5700 3064
rect 5820 3656 5828 3664
rect 5852 3856 5860 3864
rect 5900 3856 5908 3864
rect 5932 3936 5940 3944
rect 5996 4336 6004 4344
rect 6012 4316 6020 4324
rect 5996 4296 6004 4304
rect 6012 4276 6020 4284
rect 6044 4616 6052 4624
rect 6108 4696 6116 4704
rect 6140 4696 6148 4704
rect 6092 4676 6100 4684
rect 6092 4596 6100 4604
rect 6092 4556 6100 4564
rect 6060 4536 6068 4544
rect 6188 4896 6196 4904
rect 6204 4876 6212 4884
rect 6188 4836 6196 4844
rect 6124 4676 6132 4684
rect 6076 4516 6084 4524
rect 6108 4516 6116 4524
rect 6060 4336 6068 4344
rect 6060 4316 6068 4324
rect 6044 4276 6052 4284
rect 6028 4256 6036 4264
rect 6060 4236 6068 4244
rect 6044 4216 6052 4224
rect 6172 4676 6180 4684
rect 6220 4816 6228 4824
rect 6204 4696 6212 4704
rect 6156 4656 6164 4664
rect 6140 4556 6148 4564
rect 6092 4496 6100 4504
rect 6124 4496 6132 4504
rect 6204 4536 6212 4544
rect 6124 4476 6132 4484
rect 6156 4476 6164 4484
rect 6108 4336 6116 4344
rect 6092 4296 6100 4304
rect 6092 4256 6100 4264
rect 6044 4156 6052 4164
rect 6012 4136 6020 4144
rect 6028 4116 6036 4124
rect 5996 4056 6004 4064
rect 5980 3996 5988 4004
rect 5980 3956 5988 3964
rect 5964 3876 5972 3884
rect 5932 3856 5940 3864
rect 5948 3856 5956 3864
rect 5980 3856 5988 3864
rect 5948 3836 5956 3844
rect 5932 3796 5940 3804
rect 5868 3756 5876 3764
rect 5884 3716 5892 3724
rect 5916 3776 5924 3784
rect 5964 3796 5972 3804
rect 5980 3796 5988 3804
rect 5964 3776 5972 3784
rect 5948 3756 5956 3764
rect 5980 3756 5988 3764
rect 5948 3676 5956 3684
rect 5852 3656 5860 3664
rect 5836 3596 5844 3604
rect 5820 3536 5828 3544
rect 5868 3636 5876 3644
rect 5932 3636 5940 3644
rect 6172 4416 6180 4424
rect 6156 4376 6164 4384
rect 6140 4316 6148 4324
rect 6188 4356 6196 4364
rect 6204 4356 6212 4364
rect 6204 4316 6212 4324
rect 6252 4976 6260 4984
rect 6252 4936 6260 4944
rect 6252 4896 6260 4904
rect 6252 4876 6260 4884
rect 6236 4616 6244 4624
rect 6252 4436 6260 4444
rect 6252 4396 6260 4404
rect 6220 4296 6228 4304
rect 6140 4276 6148 4284
rect 6108 4156 6116 4164
rect 6124 4156 6132 4164
rect 6092 4096 6100 4104
rect 6124 4096 6132 4104
rect 6060 4056 6068 4064
rect 6092 4056 6100 4064
rect 6028 3976 6036 3984
rect 6028 3956 6036 3964
rect 6076 3956 6084 3964
rect 6060 3936 6068 3944
rect 6044 3876 6052 3884
rect 6028 3856 6036 3864
rect 6012 3836 6020 3844
rect 6076 3816 6084 3824
rect 5916 3596 5924 3604
rect 5852 3516 5860 3524
rect 5836 3456 5844 3464
rect 5852 3436 5860 3444
rect 5836 3396 5844 3404
rect 5820 3336 5828 3344
rect 5820 3256 5828 3264
rect 5724 3116 5732 3124
rect 5740 3116 5748 3124
rect 5724 3096 5732 3104
rect 5740 3096 5748 3104
rect 5644 2956 5652 2964
rect 5660 2956 5668 2964
rect 5772 3076 5780 3084
rect 5756 3056 5764 3064
rect 5820 3216 5828 3224
rect 5852 3336 5860 3344
rect 5836 3196 5844 3204
rect 5820 3176 5828 3184
rect 5900 3516 5908 3524
rect 5900 3496 5908 3504
rect 5884 3416 5892 3424
rect 5948 3576 5956 3584
rect 5932 3496 5940 3504
rect 5996 3616 6004 3624
rect 6044 3756 6052 3764
rect 6028 3676 6036 3684
rect 6012 3596 6020 3604
rect 5964 3556 5972 3564
rect 5980 3556 5988 3564
rect 5932 3476 5940 3484
rect 5916 3356 5924 3364
rect 5948 3436 5956 3444
rect 5948 3376 5956 3384
rect 5884 3336 5892 3344
rect 5900 3336 5908 3344
rect 5932 3336 5940 3344
rect 5900 3316 5908 3324
rect 6076 3656 6084 3664
rect 5996 3536 6004 3544
rect 6044 3536 6052 3544
rect 5996 3496 6004 3504
rect 6060 3496 6068 3504
rect 6060 3456 6068 3464
rect 6252 4256 6260 4264
rect 6156 4236 6164 4244
rect 6236 4236 6244 4244
rect 6188 4196 6196 4204
rect 6204 4176 6212 4184
rect 6172 4156 6180 4164
rect 6172 4116 6180 4124
rect 6172 4096 6180 4104
rect 6156 4056 6164 4064
rect 6108 4016 6116 4024
rect 6140 4016 6148 4024
rect 6124 3996 6132 4004
rect 6140 3956 6148 3964
rect 6188 4056 6196 4064
rect 6188 4036 6196 4044
rect 6172 3956 6180 3964
rect 6172 3916 6180 3924
rect 6156 3876 6164 3884
rect 6124 3856 6132 3864
rect 6140 3856 6148 3864
rect 6172 3856 6180 3864
rect 6156 3836 6164 3844
rect 6124 3796 6132 3804
rect 6156 3776 6164 3784
rect 6140 3756 6148 3764
rect 6124 3716 6132 3724
rect 6108 3696 6116 3704
rect 6124 3656 6132 3664
rect 6156 3716 6164 3724
rect 6188 3796 6196 3804
rect 6188 3776 6196 3784
rect 6188 3736 6196 3744
rect 6172 3696 6180 3704
rect 6092 3636 6100 3644
rect 6124 3636 6132 3644
rect 6140 3636 6148 3644
rect 6108 3616 6116 3624
rect 6108 3516 6116 3524
rect 6140 3576 6148 3584
rect 6188 3636 6196 3644
rect 6172 3516 6180 3524
rect 6124 3496 6132 3504
rect 6188 3496 6196 3504
rect 6172 3476 6180 3484
rect 5980 3436 5988 3444
rect 6076 3436 6084 3444
rect 6108 3436 6116 3444
rect 5964 3336 5972 3344
rect 6028 3416 6036 3424
rect 5996 3376 6004 3384
rect 5900 3276 5908 3284
rect 5916 3276 5924 3284
rect 5836 3136 5844 3144
rect 5868 3136 5876 3144
rect 5820 3096 5828 3104
rect 5804 3076 5812 3084
rect 5900 3236 5908 3244
rect 5916 3216 5924 3224
rect 5916 3156 5924 3164
rect 5900 3116 5908 3124
rect 5868 3096 5876 3104
rect 5756 3016 5764 3024
rect 5788 3016 5796 3024
rect 5756 2956 5764 2964
rect 5548 2816 5556 2824
rect 5532 2776 5540 2784
rect 5468 2756 5476 2764
rect 5500 2756 5508 2764
rect 5516 2756 5524 2764
rect 5836 3036 5844 3044
rect 5884 3036 5892 3044
rect 5836 3016 5844 3024
rect 5804 2976 5812 2984
rect 5820 2976 5828 2984
rect 5868 2976 5876 2984
rect 5788 2956 5796 2964
rect 5804 2956 5812 2964
rect 5676 2936 5684 2944
rect 5724 2936 5732 2944
rect 5708 2896 5716 2904
rect 5612 2836 5620 2844
rect 5596 2816 5604 2824
rect 5564 2716 5572 2724
rect 5564 2696 5572 2704
rect 5644 2696 5652 2704
rect 5660 2696 5668 2704
rect 5532 2676 5540 2684
rect 5580 2676 5588 2684
rect 5628 2676 5636 2684
rect 5596 2656 5604 2664
rect 5612 2656 5620 2664
rect 5596 2636 5604 2644
rect 5692 2776 5700 2784
rect 5724 2836 5732 2844
rect 5756 2896 5764 2904
rect 5788 2896 5796 2904
rect 5804 2896 5812 2904
rect 5756 2836 5764 2844
rect 5756 2816 5764 2824
rect 5772 2816 5780 2824
rect 5804 2816 5812 2824
rect 5740 2776 5748 2784
rect 5900 2956 5908 2964
rect 5788 2776 5796 2784
rect 5820 2776 5828 2784
rect 5756 2736 5764 2744
rect 5772 2736 5780 2744
rect 5708 2716 5716 2724
rect 5724 2716 5732 2724
rect 5692 2696 5700 2704
rect 5692 2676 5700 2684
rect 5756 2696 5764 2704
rect 5772 2676 5780 2684
rect 5740 2656 5748 2664
rect 5756 2656 5764 2664
rect 5660 2636 5668 2644
rect 5676 2636 5684 2644
rect 5724 2636 5732 2644
rect 5468 2536 5476 2544
rect 5468 2476 5476 2484
rect 5452 2376 5460 2384
rect 5324 2336 5332 2344
rect 5404 2336 5412 2344
rect 5468 2316 5476 2324
rect 5324 2296 5332 2304
rect 5356 2296 5364 2304
rect 5180 2276 5188 2284
rect 5292 2276 5300 2284
rect 5308 2276 5316 2284
rect 5436 2276 5444 2284
rect 5148 2256 5156 2264
rect 5276 2256 5284 2264
rect 5036 2156 5044 2164
rect 5068 2176 5076 2184
rect 5468 2256 5476 2264
rect 5324 2236 5332 2244
rect 5244 2216 5252 2224
rect 5148 2196 5156 2204
rect 5212 2196 5220 2204
rect 5100 2176 5108 2184
rect 5132 2176 5140 2184
rect 5132 2156 5140 2164
rect 5148 2136 5156 2144
rect 5004 2116 5012 2124
rect 5052 2116 5060 2124
rect 5068 2116 5076 2124
rect 5132 2116 5140 2124
rect 5228 2136 5236 2144
rect 5324 2176 5332 2184
rect 5388 2176 5396 2184
rect 5340 2156 5348 2164
rect 5292 2136 5300 2144
rect 5548 2616 5556 2624
rect 5564 2536 5572 2544
rect 5580 2536 5588 2544
rect 5708 2536 5716 2544
rect 5516 2516 5524 2524
rect 5532 2516 5540 2524
rect 5596 2516 5604 2524
rect 5660 2516 5668 2524
rect 5500 2476 5508 2484
rect 5516 2476 5524 2484
rect 5548 2456 5556 2464
rect 5532 2416 5540 2424
rect 5580 2416 5588 2424
rect 5548 2356 5556 2364
rect 5660 2376 5668 2384
rect 5564 2316 5572 2324
rect 5628 2316 5636 2324
rect 5900 2916 5908 2924
rect 5868 2856 5876 2864
rect 5852 2836 5860 2844
rect 5868 2836 5876 2844
rect 5852 2816 5860 2824
rect 5804 2716 5812 2724
rect 5836 2716 5844 2724
rect 5788 2616 5796 2624
rect 5820 2696 5828 2704
rect 5820 2676 5828 2684
rect 5756 2576 5764 2584
rect 5788 2556 5796 2564
rect 5740 2496 5748 2504
rect 5772 2456 5780 2464
rect 5788 2456 5796 2464
rect 5500 2276 5508 2284
rect 5660 2296 5668 2304
rect 5724 2296 5732 2304
rect 5692 2276 5700 2284
rect 5548 2256 5556 2264
rect 5596 2256 5604 2264
rect 5868 2736 5876 2744
rect 5980 3296 5988 3304
rect 6012 3336 6020 3344
rect 5964 3256 5972 3264
rect 5996 3276 6004 3284
rect 6012 3276 6020 3284
rect 6012 3176 6020 3184
rect 5980 3156 5988 3164
rect 5964 3096 5972 3104
rect 5932 2976 5940 2984
rect 5948 2976 5956 2984
rect 6012 3136 6020 3144
rect 6060 3396 6068 3404
rect 6140 3396 6148 3404
rect 6188 3456 6196 3464
rect 6172 3356 6180 3364
rect 6220 4076 6228 4084
rect 6236 3996 6244 4004
rect 6220 3896 6228 3904
rect 6220 3776 6228 3784
rect 6220 3756 6228 3764
rect 6220 3736 6228 3744
rect 6236 3736 6244 3744
rect 6236 3716 6244 3724
rect 6220 3696 6228 3704
rect 6220 3656 6228 3664
rect 6220 3596 6228 3604
rect 6220 3536 6228 3544
rect 6220 3516 6228 3524
rect 6220 3476 6228 3484
rect 6220 3456 6228 3464
rect 6204 3396 6212 3404
rect 6220 3376 6228 3384
rect 6220 3356 6228 3364
rect 6124 3316 6132 3324
rect 6060 3276 6068 3284
rect 6028 3116 6036 3124
rect 6028 3076 6036 3084
rect 6124 3216 6132 3224
rect 6076 3116 6084 3124
rect 6092 3096 6100 3104
rect 6028 3036 6036 3044
rect 6060 3036 6068 3044
rect 5996 2976 6004 2984
rect 5932 2956 5940 2964
rect 5948 2956 5956 2964
rect 5980 2956 5988 2964
rect 5980 2936 5988 2944
rect 5948 2916 5956 2924
rect 5964 2916 5972 2924
rect 6012 2936 6020 2944
rect 5948 2876 5956 2884
rect 5964 2836 5972 2844
rect 5980 2836 5988 2844
rect 5948 2816 5956 2824
rect 5900 2696 5908 2704
rect 5884 2676 5892 2684
rect 5900 2676 5908 2684
rect 5852 2656 5860 2664
rect 5836 2636 5844 2644
rect 5836 2616 5844 2624
rect 5852 2616 5860 2624
rect 5916 2616 5924 2624
rect 5836 2556 5844 2564
rect 5852 2536 5860 2544
rect 5836 2516 5844 2524
rect 5804 2356 5812 2364
rect 5644 2216 5652 2224
rect 5708 2216 5716 2224
rect 5740 2216 5748 2224
rect 5404 2156 5412 2164
rect 5484 2156 5492 2164
rect 5628 2156 5636 2164
rect 5356 2136 5364 2144
rect 5244 2116 5252 2124
rect 5276 2116 5284 2124
rect 5148 2076 5156 2084
rect 5308 2076 5316 2084
rect 5292 2056 5300 2064
rect 5628 2136 5636 2144
rect 5436 2116 5444 2124
rect 5516 2116 5524 2124
rect 5564 2116 5572 2124
rect 5388 2096 5396 2104
rect 5356 2036 5364 2044
rect 5372 2036 5380 2044
rect 4956 2016 4964 2024
rect 4988 2016 4996 2024
rect 4940 1996 4948 2004
rect 4940 1956 4948 1964
rect 4908 1916 4916 1924
rect 5260 1976 5268 1984
rect 5148 1916 5156 1924
rect 5180 1916 5188 1924
rect 4956 1896 4964 1904
rect 5020 1896 5028 1904
rect 5132 1896 5140 1904
rect 4828 1856 4836 1864
rect 4860 1856 4868 1864
rect 5036 1856 5044 1864
rect 4828 1796 4836 1804
rect 4940 1796 4948 1804
rect 4876 1776 4884 1784
rect 4988 1776 4996 1784
rect 5148 1856 5156 1864
rect 5180 1856 5188 1864
rect 5244 1876 5252 1884
rect 5228 1856 5236 1864
rect 5196 1836 5204 1844
rect 5212 1836 5220 1844
rect 5484 2056 5492 2064
rect 5580 2076 5588 2084
rect 5756 2196 5764 2204
rect 5804 2236 5812 2244
rect 5660 2116 5668 2124
rect 5724 2116 5732 2124
rect 5676 2096 5684 2104
rect 5708 2096 5716 2104
rect 5772 2096 5780 2104
rect 5724 2076 5732 2084
rect 5612 2056 5620 2064
rect 5644 2056 5652 2064
rect 5468 2036 5476 2044
rect 5500 2036 5508 2044
rect 5532 2036 5540 2044
rect 5372 1956 5380 1964
rect 5420 1956 5428 1964
rect 5276 1856 5284 1864
rect 5356 1856 5364 1864
rect 5292 1836 5300 1844
rect 5324 1836 5332 1844
rect 5500 2016 5508 2024
rect 5532 2016 5540 2024
rect 5468 1956 5476 1964
rect 5484 1956 5492 1964
rect 5452 1916 5460 1924
rect 5484 1916 5492 1924
rect 5548 1936 5556 1944
rect 5580 1916 5588 1924
rect 5388 1876 5396 1884
rect 5532 1876 5540 1884
rect 5420 1856 5428 1864
rect 5276 1816 5284 1824
rect 5372 1816 5380 1824
rect 5820 2216 5828 2224
rect 5804 2036 5812 2044
rect 5740 2016 5748 2024
rect 5772 2016 5780 2024
rect 5660 1916 5668 1924
rect 5596 1856 5604 1864
rect 5340 1776 5348 1784
rect 4924 1756 4932 1764
rect 4972 1756 4980 1764
rect 5068 1756 5076 1764
rect 5260 1756 5268 1764
rect 5292 1756 5300 1764
rect 5484 1756 5492 1764
rect 5564 1756 5572 1764
rect 4796 1736 4804 1744
rect 4748 1656 4756 1664
rect 4812 1596 4820 1604
rect 4876 1716 4884 1724
rect 4892 1716 4900 1724
rect 5068 1736 5076 1744
rect 5132 1736 5140 1744
rect 5308 1736 5316 1744
rect 4876 1696 4884 1704
rect 4828 1556 4836 1564
rect 4764 1516 4772 1524
rect 4828 1516 4836 1524
rect 4732 1496 4740 1504
rect 4748 1496 4756 1504
rect 4716 1476 4724 1484
rect 4812 1496 4820 1504
rect 4860 1496 4868 1504
rect 4876 1496 4884 1504
rect 4636 1456 4644 1464
rect 4668 1456 4676 1464
rect 4556 1436 4564 1444
rect 4796 1436 4804 1444
rect 4844 1436 4852 1444
rect 4540 1416 4548 1424
rect 4780 1416 4788 1424
rect 4492 1356 4500 1364
rect 4764 1336 4772 1344
rect 4556 1316 4564 1324
rect 4492 1296 4500 1304
rect 4524 1276 4532 1284
rect 4476 1256 4484 1264
rect 4444 1236 4452 1244
rect 4396 1156 4404 1164
rect 4348 1136 4356 1144
rect 3980 1076 3988 1084
rect 4108 1096 4116 1104
rect 3932 1056 3940 1064
rect 3996 1056 4004 1064
rect 4060 1056 4068 1064
rect 4076 1056 4084 1064
rect 3884 1016 3892 1024
rect 3820 976 3828 984
rect 3836 976 3844 984
rect 3868 976 3876 984
rect 3852 956 3860 964
rect 3708 936 3716 944
rect 3804 936 3812 944
rect 3868 936 3876 944
rect 3404 916 3412 924
rect 3516 916 3524 924
rect 3660 916 3668 924
rect 3436 896 3444 904
rect 3388 816 3396 824
rect 3404 816 3412 824
rect 3388 756 3396 764
rect 3356 716 3364 724
rect 3292 696 3300 704
rect 3356 696 3364 704
rect 3500 856 3508 864
rect 3452 836 3460 844
rect 3404 716 3412 724
rect 3500 736 3508 744
rect 3276 636 3284 644
rect 3388 636 3396 644
rect 3180 616 3188 624
rect 3118 606 3126 614
rect 3132 606 3140 614
rect 3146 606 3154 614
rect 3148 576 3156 584
rect 3116 536 3124 544
rect 3244 556 3252 564
rect 3276 556 3284 564
rect 3180 536 3188 544
rect 3244 536 3252 544
rect 3164 496 3172 504
rect 3164 476 3172 484
rect 3212 496 3220 504
rect 3404 616 3412 624
rect 3468 696 3476 704
rect 3548 696 3556 704
rect 3564 696 3572 704
rect 3788 916 3796 924
rect 3644 896 3652 904
rect 3676 896 3684 904
rect 3804 896 3812 904
rect 3740 876 3748 884
rect 3772 876 3780 884
rect 3676 736 3684 744
rect 3708 736 3716 744
rect 3724 736 3732 744
rect 3740 716 3748 724
rect 3644 696 3652 704
rect 3660 696 3668 704
rect 3724 696 3732 704
rect 3772 696 3780 704
rect 3596 676 3604 684
rect 3612 676 3620 684
rect 3452 656 3460 664
rect 3420 556 3428 564
rect 3292 516 3300 524
rect 3292 496 3300 504
rect 3372 496 3380 504
rect 3260 456 3268 464
rect 3308 456 3316 464
rect 3356 376 3364 384
rect 3212 316 3220 324
rect 3324 316 3332 324
rect 3372 316 3380 324
rect 3420 316 3428 324
rect 3148 276 3156 284
rect 3468 496 3476 504
rect 3516 656 3524 664
rect 3580 656 3588 664
rect 3660 656 3668 664
rect 3500 636 3508 644
rect 3532 636 3540 644
rect 3580 636 3588 644
rect 3708 616 3716 624
rect 3804 816 3812 824
rect 3836 756 3844 764
rect 3820 696 3828 704
rect 3804 656 3812 664
rect 3852 656 3860 664
rect 3788 576 3796 584
rect 3500 556 3508 564
rect 3612 556 3620 564
rect 3724 556 3732 564
rect 3836 556 3844 564
rect 3708 536 3716 544
rect 3820 536 3828 544
rect 3516 496 3524 504
rect 4028 976 4036 984
rect 4060 976 4068 984
rect 3948 956 3956 964
rect 4092 956 4100 964
rect 3916 936 3924 944
rect 3932 916 3940 924
rect 4044 936 4052 944
rect 3996 916 4004 924
rect 4028 916 4036 924
rect 3900 896 3908 904
rect 3916 876 3924 884
rect 3980 876 3988 884
rect 3932 856 3940 864
rect 3900 756 3908 764
rect 3916 736 3924 744
rect 3916 696 3924 704
rect 3964 736 3972 744
rect 3948 696 3956 704
rect 4012 736 4020 744
rect 3980 696 3988 704
rect 3996 696 4004 704
rect 4188 1116 4196 1124
rect 4380 1116 4388 1124
rect 4156 996 4164 1004
rect 4252 1096 4260 1104
rect 4412 1096 4420 1104
rect 4220 1076 4228 1084
rect 4284 1076 4292 1084
rect 4252 1056 4260 1064
rect 4268 1056 4276 1064
rect 4300 1056 4308 1064
rect 4300 1036 4308 1044
rect 4364 1016 4372 1024
rect 4412 1016 4420 1024
rect 4492 1116 4500 1124
rect 4460 1096 4468 1104
rect 4556 1096 4564 1104
rect 4588 1076 4596 1084
rect 4476 1036 4484 1044
rect 4796 1316 4804 1324
rect 4636 1296 4644 1304
rect 4764 1296 4772 1304
rect 4828 1336 4836 1344
rect 4716 1276 4724 1284
rect 4638 1206 4646 1214
rect 4652 1206 4660 1214
rect 4666 1206 4674 1214
rect 4908 1696 4916 1704
rect 4988 1716 4996 1724
rect 5004 1716 5012 1724
rect 5036 1716 5044 1724
rect 4956 1656 4964 1664
rect 5084 1656 5092 1664
rect 4988 1636 4996 1644
rect 5308 1716 5316 1724
rect 5388 1736 5396 1744
rect 5404 1716 5412 1724
rect 5420 1716 5428 1724
rect 5468 1716 5476 1724
rect 5356 1696 5364 1704
rect 5372 1696 5380 1704
rect 5516 1740 5524 1744
rect 5516 1736 5524 1740
rect 5500 1716 5508 1724
rect 5596 1716 5604 1724
rect 5596 1696 5604 1704
rect 5452 1636 5460 1644
rect 5148 1616 5156 1624
rect 5260 1616 5268 1624
rect 5468 1616 5476 1624
rect 5036 1596 5044 1604
rect 4956 1576 4964 1584
rect 4924 1556 4932 1564
rect 4908 1536 4916 1544
rect 4956 1536 4964 1544
rect 4972 1516 4980 1524
rect 5020 1516 5028 1524
rect 4924 1496 4932 1504
rect 4940 1496 4948 1504
rect 5004 1496 5012 1504
rect 4892 1476 4900 1484
rect 4972 1476 4980 1484
rect 5004 1456 5012 1464
rect 4988 1436 4996 1444
rect 4876 1356 4884 1364
rect 4940 1356 4948 1364
rect 5308 1556 5316 1564
rect 5356 1556 5364 1564
rect 5100 1536 5108 1544
rect 5292 1536 5300 1544
rect 5068 1516 5076 1524
rect 5132 1516 5140 1524
rect 5164 1516 5172 1524
rect 5052 1496 5060 1504
rect 5100 1496 5108 1504
rect 5052 1456 5060 1464
rect 5340 1536 5348 1544
rect 5196 1496 5204 1504
rect 5356 1516 5364 1524
rect 5436 1516 5444 1524
rect 5436 1496 5444 1504
rect 5564 1496 5572 1504
rect 5420 1476 5428 1484
rect 5276 1456 5284 1464
rect 5324 1456 5332 1464
rect 5388 1456 5396 1464
rect 5404 1456 5412 1464
rect 5084 1416 5092 1424
rect 5180 1416 5188 1424
rect 5132 1396 5140 1404
rect 5052 1336 5060 1344
rect 5196 1356 5204 1364
rect 5260 1356 5268 1364
rect 5212 1336 5220 1344
rect 5244 1336 5252 1344
rect 4892 1316 4900 1324
rect 5004 1316 5012 1324
rect 5020 1316 5028 1324
rect 5100 1316 5108 1324
rect 5084 1296 5092 1304
rect 5052 1256 5060 1264
rect 4860 1176 4868 1184
rect 4636 1116 4644 1124
rect 4716 1116 4724 1124
rect 4908 1116 4916 1124
rect 4780 1096 4788 1104
rect 4844 1096 4852 1104
rect 4828 1076 4836 1084
rect 4732 1056 4740 1064
rect 4940 1156 4948 1164
rect 4956 1116 4964 1124
rect 4892 1076 4900 1084
rect 4924 1076 4932 1084
rect 4988 1156 4996 1164
rect 5052 1096 5060 1104
rect 5484 1476 5492 1484
rect 5532 1476 5540 1484
rect 5468 1436 5476 1444
rect 5308 1316 5316 1324
rect 5164 1296 5172 1304
rect 5436 1336 5444 1344
rect 5660 1896 5668 1904
rect 5708 1956 5716 1964
rect 5692 1936 5700 1944
rect 5724 1896 5732 1904
rect 5708 1876 5716 1884
rect 5772 1876 5780 1884
rect 5900 2556 5908 2564
rect 5948 2736 5956 2744
rect 5964 2676 5972 2684
rect 5948 2596 5956 2604
rect 6012 2756 6020 2764
rect 6012 2736 6020 2744
rect 6060 3016 6068 3024
rect 6156 3116 6164 3124
rect 6156 3076 6164 3084
rect 6188 3316 6196 3324
rect 6236 3316 6244 3324
rect 6236 3116 6244 3124
rect 6156 3056 6164 3064
rect 6172 3056 6180 3064
rect 6204 3056 6212 3064
rect 6124 2976 6132 2984
rect 6092 2956 6100 2964
rect 6076 2916 6084 2924
rect 6060 2876 6068 2884
rect 6108 2936 6116 2944
rect 6108 2916 6116 2924
rect 6060 2856 6068 2864
rect 6092 2856 6100 2864
rect 6044 2756 6052 2764
rect 6012 2696 6020 2704
rect 6028 2696 6036 2704
rect 6012 2676 6020 2684
rect 6028 2676 6036 2684
rect 6044 2676 6052 2684
rect 5996 2616 6004 2624
rect 6028 2636 6036 2644
rect 5980 2576 5988 2584
rect 5996 2576 6004 2584
rect 6012 2576 6020 2584
rect 5884 2476 5892 2484
rect 5884 2456 5892 2464
rect 5916 2536 5924 2544
rect 5932 2516 5940 2524
rect 5996 2516 6004 2524
rect 6028 2516 6036 2524
rect 6044 2516 6052 2524
rect 5932 2496 5940 2504
rect 5980 2496 5988 2504
rect 5916 2476 5924 2484
rect 5948 2476 5956 2484
rect 5932 2456 5940 2464
rect 5852 2356 5860 2364
rect 5868 2356 5876 2364
rect 5900 2396 5908 2404
rect 5900 2376 5908 2384
rect 5868 2276 5876 2284
rect 5852 2236 5860 2244
rect 5884 2236 5892 2244
rect 5836 2116 5844 2124
rect 5868 2096 5876 2104
rect 5868 2076 5876 2084
rect 5884 2076 5892 2084
rect 5820 1856 5828 1864
rect 5788 1836 5796 1844
rect 5628 1776 5636 1784
rect 5708 1776 5716 1784
rect 5644 1716 5652 1724
rect 5676 1696 5684 1704
rect 5740 1716 5748 1724
rect 5820 1796 5828 1804
rect 5852 1956 5860 1964
rect 5916 2296 5924 2304
rect 5932 2296 5940 2304
rect 5900 1996 5908 2004
rect 5884 1916 5892 1924
rect 5932 2236 5940 2244
rect 5948 2176 5956 2184
rect 5948 2156 5956 2164
rect 5932 2116 5940 2124
rect 5996 2396 6004 2404
rect 5996 2376 6004 2384
rect 6076 2716 6084 2724
rect 6092 2696 6100 2704
rect 6076 2636 6084 2644
rect 6076 2596 6084 2604
rect 6124 2896 6132 2904
rect 6124 2876 6132 2884
rect 6124 2796 6132 2804
rect 6124 2696 6132 2704
rect 6156 2916 6164 2924
rect 6188 2916 6196 2924
rect 6172 2816 6180 2824
rect 6156 2716 6164 2724
rect 6172 2716 6180 2724
rect 6124 2676 6132 2684
rect 6140 2676 6148 2684
rect 6172 2676 6180 2684
rect 6092 2556 6100 2564
rect 6108 2556 6116 2564
rect 6108 2536 6116 2544
rect 6092 2456 6100 2464
rect 6076 2416 6084 2424
rect 6060 2396 6068 2404
rect 6012 2356 6020 2364
rect 6028 2356 6036 2364
rect 5996 2336 6004 2344
rect 5980 2236 5988 2244
rect 5980 2216 5988 2224
rect 5980 2136 5988 2144
rect 5964 1976 5972 1984
rect 5932 1956 5940 1964
rect 5948 1956 5956 1964
rect 5932 1936 5940 1944
rect 6012 2276 6020 2284
rect 6044 2316 6052 2324
rect 6028 2196 6036 2204
rect 6060 2276 6068 2284
rect 6076 2276 6084 2284
rect 6060 2236 6068 2244
rect 6012 2136 6020 2144
rect 6044 2136 6052 2144
rect 6012 2116 6020 2124
rect 6028 2096 6036 2104
rect 6076 2196 6084 2204
rect 6108 2336 6116 2344
rect 6108 2316 6116 2324
rect 6140 2656 6148 2664
rect 6140 2636 6148 2644
rect 6156 2616 6164 2624
rect 6156 2516 6164 2524
rect 6140 2416 6148 2424
rect 6156 2376 6164 2384
rect 6236 3036 6244 3044
rect 6236 2936 6244 2944
rect 6220 2836 6228 2844
rect 6220 2816 6228 2824
rect 6236 2776 6244 2784
rect 6204 2736 6212 2744
rect 6220 2716 6228 2724
rect 6204 2696 6212 2704
rect 6188 2616 6196 2624
rect 6188 2576 6196 2584
rect 6204 2476 6212 2484
rect 6188 2356 6196 2364
rect 6172 2296 6180 2304
rect 6124 2276 6132 2284
rect 6140 2236 6148 2244
rect 6188 2236 6196 2244
rect 6140 2196 6148 2204
rect 6108 2176 6116 2184
rect 6044 2076 6052 2084
rect 5996 1936 6004 1944
rect 5868 1896 5876 1904
rect 5868 1876 5876 1884
rect 5932 1896 5940 1904
rect 5916 1876 5924 1884
rect 5884 1856 5892 1864
rect 5900 1856 5908 1864
rect 5916 1816 5924 1824
rect 5724 1696 5732 1704
rect 5804 1696 5812 1704
rect 5740 1616 5748 1624
rect 5692 1536 5700 1544
rect 5724 1516 5732 1524
rect 5692 1496 5700 1504
rect 5580 1456 5588 1464
rect 5612 1456 5620 1464
rect 5580 1436 5588 1444
rect 5580 1396 5588 1404
rect 5580 1316 5588 1324
rect 5628 1316 5636 1324
rect 5884 1776 5892 1784
rect 5932 1796 5940 1804
rect 5980 1916 5988 1924
rect 5980 1876 5988 1884
rect 5964 1836 5972 1844
rect 5996 1776 6004 1784
rect 5948 1756 5956 1764
rect 5948 1736 5956 1744
rect 5948 1716 5956 1724
rect 5836 1676 5844 1684
rect 5884 1696 5892 1704
rect 5852 1656 5860 1664
rect 5836 1536 5844 1544
rect 5788 1516 5796 1524
rect 5820 1516 5828 1524
rect 5980 1696 5988 1704
rect 5948 1576 5956 1584
rect 5932 1536 5940 1544
rect 5740 1496 5748 1504
rect 5820 1496 5828 1504
rect 5868 1496 5876 1504
rect 5788 1476 5796 1484
rect 5884 1476 5892 1484
rect 5708 1436 5716 1444
rect 5772 1436 5780 1444
rect 5756 1376 5764 1384
rect 5756 1356 5764 1364
rect 5692 1336 5700 1344
rect 5756 1336 5764 1344
rect 5340 1296 5348 1304
rect 5420 1296 5428 1304
rect 5596 1296 5604 1304
rect 5660 1316 5668 1324
rect 5756 1316 5764 1324
rect 5644 1296 5652 1304
rect 5500 1276 5508 1284
rect 5564 1276 5572 1284
rect 5612 1276 5620 1284
rect 5244 1236 5252 1244
rect 5292 1236 5300 1244
rect 5148 1176 5156 1184
rect 5244 1176 5252 1184
rect 5180 1156 5188 1164
rect 5260 1136 5268 1144
rect 5132 1116 5140 1124
rect 5228 1116 5236 1124
rect 5004 1076 5012 1084
rect 5228 1096 5236 1104
rect 4972 1056 4980 1064
rect 5132 1056 5140 1064
rect 4748 1036 4756 1044
rect 4860 1036 4868 1044
rect 4988 1036 4996 1044
rect 4604 996 4612 1004
rect 4444 976 4452 984
rect 4540 976 4548 984
rect 4588 976 4596 984
rect 4876 976 4884 984
rect 4908 976 4916 984
rect 4220 956 4228 964
rect 4396 956 4404 964
rect 4428 956 4436 964
rect 4460 956 4468 964
rect 4524 956 4532 964
rect 4332 936 4340 944
rect 4380 936 4388 944
rect 4428 936 4436 944
rect 4476 936 4484 944
rect 4524 936 4532 944
rect 4556 936 4564 944
rect 4572 936 4580 944
rect 4700 956 4708 964
rect 4748 956 4756 964
rect 4796 956 4804 964
rect 4844 936 4852 944
rect 4892 936 4900 944
rect 4956 936 4964 944
rect 4156 696 4164 704
rect 4684 916 4692 924
rect 4732 916 4740 924
rect 4908 916 4916 924
rect 4236 896 4244 904
rect 4348 896 4356 904
rect 4460 896 4468 904
rect 4508 896 4516 904
rect 4796 896 4804 904
rect 4860 896 4868 904
rect 4012 676 4020 684
rect 4028 676 4036 684
rect 4140 676 4148 684
rect 4172 676 4180 684
rect 3932 636 3940 644
rect 3948 596 3956 604
rect 3916 556 3924 564
rect 3932 556 3940 564
rect 3868 536 3876 544
rect 3980 556 3988 564
rect 3964 536 3972 544
rect 3804 496 3812 504
rect 4188 656 4196 664
rect 4092 636 4100 644
rect 4044 576 4052 584
rect 4012 536 4020 544
rect 3868 476 3876 484
rect 3900 476 3908 484
rect 3948 476 3956 484
rect 4076 536 4084 544
rect 3852 456 3860 464
rect 3884 456 3892 464
rect 3692 436 3700 444
rect 3676 416 3684 424
rect 3484 336 3492 344
rect 3532 336 3540 344
rect 3660 336 3668 344
rect 3388 296 3396 304
rect 3452 296 3460 304
rect 3500 296 3508 304
rect 3228 276 3236 284
rect 3340 276 3348 284
rect 3484 276 3492 284
rect 3580 316 3588 324
rect 3660 296 3668 304
rect 3516 256 3524 264
rect 3180 236 3188 244
rect 3292 236 3300 244
rect 3118 206 3126 214
rect 3132 206 3140 214
rect 3146 206 3154 214
rect 3084 196 3092 204
rect 3532 196 3540 204
rect 3596 196 3604 204
rect 3612 196 3620 204
rect 2476 176 2484 184
rect 2604 136 2612 144
rect 2652 136 2660 144
rect 2748 156 2756 164
rect 2812 156 2820 164
rect 2892 156 2900 164
rect 2924 156 2932 164
rect 3196 156 3204 164
rect 3308 156 3316 164
rect 3500 156 3508 164
rect 2524 116 2532 124
rect 2508 16 2516 24
rect 2620 116 2628 124
rect 2668 116 2676 124
rect 2700 116 2708 124
rect 2716 116 2724 124
rect 2796 116 2804 124
rect 2764 96 2772 104
rect 2780 96 2788 104
rect 2780 56 2788 64
rect 2908 116 2916 124
rect 2876 96 2884 104
rect 3052 136 3060 144
rect 3116 136 3124 144
rect 3452 136 3460 144
rect 2972 96 2980 104
rect 3068 116 3076 124
rect 3212 116 3220 124
rect 3052 96 3060 104
rect 3180 96 3188 104
rect 3308 116 3316 124
rect 3340 116 3348 124
rect 3452 116 3460 124
rect 3260 96 3268 104
rect 3436 56 3444 64
rect 3692 396 3700 404
rect 3996 436 4004 444
rect 3900 396 3908 404
rect 4012 396 4020 404
rect 4028 396 4036 404
rect 3788 356 3796 364
rect 3836 356 3844 364
rect 3692 296 3700 304
rect 3868 296 3876 304
rect 3708 276 3716 284
rect 3932 376 3940 384
rect 3980 376 3988 384
rect 3948 336 3956 344
rect 3964 316 3972 324
rect 4044 356 4052 364
rect 3996 316 4004 324
rect 4028 316 4036 324
rect 4108 576 4116 584
rect 4172 576 4180 584
rect 4124 536 4132 544
rect 4156 456 4164 464
rect 4188 536 4196 544
rect 4732 876 4740 884
rect 4556 736 4564 744
rect 4252 716 4260 724
rect 4300 716 4308 724
rect 4364 696 4372 704
rect 4332 676 4340 684
rect 4236 576 4244 584
rect 4268 576 4276 584
rect 4284 556 4292 564
rect 4204 516 4212 524
rect 4188 476 4196 484
rect 4140 376 4148 384
rect 4124 356 4132 364
rect 4108 316 4116 324
rect 4140 316 4148 324
rect 3948 276 3956 284
rect 3996 276 4004 284
rect 4028 276 4036 284
rect 4092 276 4100 284
rect 3756 256 3764 264
rect 3804 256 3812 264
rect 4012 256 4020 264
rect 3644 156 3652 164
rect 3644 136 3652 144
rect 3692 136 3700 144
rect 3772 216 3780 224
rect 4140 236 4148 244
rect 3900 196 3908 204
rect 4012 196 4020 204
rect 4108 196 4116 204
rect 4220 416 4228 424
rect 4252 416 4260 424
rect 4236 396 4244 404
rect 4444 716 4452 724
rect 4476 716 4484 724
rect 4572 716 4580 724
rect 4444 696 4452 704
rect 4524 696 4532 704
rect 4556 696 4564 704
rect 4396 676 4404 684
rect 4380 636 4388 644
rect 4396 636 4404 644
rect 4476 576 4484 584
rect 4332 556 4340 564
rect 4412 556 4420 564
rect 4460 556 4468 564
rect 4300 516 4308 524
rect 4364 516 4372 524
rect 4348 496 4356 504
rect 4332 476 4340 484
rect 4444 516 4452 524
rect 4460 516 4468 524
rect 4508 516 4516 524
rect 4492 496 4500 504
rect 4476 476 4484 484
rect 4380 436 4388 444
rect 4428 436 4436 444
rect 4460 436 4468 444
rect 4364 416 4372 424
rect 4364 336 4372 344
rect 4316 316 4324 324
rect 4348 316 4356 324
rect 4428 316 4436 324
rect 4268 276 4276 284
rect 4638 806 4646 814
rect 4652 806 4660 814
rect 4666 806 4674 814
rect 4924 876 4932 884
rect 4812 756 4820 764
rect 4700 736 4708 744
rect 4748 736 4756 744
rect 4780 736 4788 744
rect 5036 996 5044 1004
rect 5052 976 5060 984
rect 5020 956 5028 964
rect 5052 936 5060 944
rect 5004 916 5012 924
rect 5132 1016 5140 1024
rect 5084 976 5092 984
rect 5116 976 5124 984
rect 5068 916 5076 924
rect 5116 956 5124 964
rect 5276 1096 5284 1104
rect 5692 1156 5700 1164
rect 5340 1136 5348 1144
rect 5452 1136 5460 1144
rect 5596 1136 5604 1144
rect 5324 1076 5332 1084
rect 5276 1056 5284 1064
rect 5196 1036 5204 1044
rect 5244 1016 5252 1024
rect 5372 1096 5380 1104
rect 5404 1076 5412 1084
rect 5292 1036 5300 1044
rect 5356 1036 5364 1044
rect 5404 1036 5412 1044
rect 5516 1076 5524 1084
rect 5580 1076 5588 1084
rect 5660 1056 5668 1064
rect 5484 1016 5492 1024
rect 5436 996 5444 1004
rect 5484 996 5492 1004
rect 5180 976 5188 984
rect 5292 976 5300 984
rect 5308 976 5316 984
rect 5404 976 5412 984
rect 5148 956 5156 964
rect 5148 936 5156 944
rect 5100 896 5108 904
rect 5100 876 5108 884
rect 4972 756 4980 764
rect 4972 736 4980 744
rect 5196 936 5204 944
rect 5244 936 5252 944
rect 5180 876 5188 884
rect 5228 916 5236 924
rect 5340 916 5348 924
rect 5388 916 5396 924
rect 5452 916 5460 924
rect 5500 916 5508 924
rect 5212 896 5220 904
rect 5356 896 5364 904
rect 5388 876 5396 884
rect 5468 856 5476 864
rect 5196 836 5204 844
rect 5292 736 5300 744
rect 5324 736 5332 744
rect 5340 736 5348 744
rect 4668 716 4676 724
rect 4844 716 4852 724
rect 5004 716 5012 724
rect 5084 716 5092 724
rect 5164 716 5172 724
rect 5356 716 5364 724
rect 4604 696 4612 704
rect 4684 696 4692 704
rect 4732 696 4740 704
rect 4796 696 4804 704
rect 4908 696 4916 704
rect 4540 676 4548 684
rect 4540 656 4548 664
rect 4540 616 4548 624
rect 4556 576 4564 584
rect 4540 536 4548 544
rect 4796 676 4804 684
rect 4588 656 4596 664
rect 4732 656 4740 664
rect 4876 656 4884 664
rect 4956 656 4964 664
rect 4716 616 4724 624
rect 4796 616 4804 624
rect 4764 576 4772 584
rect 4780 576 4788 584
rect 4620 556 4628 564
rect 4636 536 4644 544
rect 4764 536 4772 544
rect 4588 496 4596 504
rect 4748 496 4756 504
rect 4812 536 4820 544
rect 4844 536 4852 544
rect 4860 496 4868 504
rect 4524 416 4532 424
rect 4540 416 4548 424
rect 4572 416 4580 424
rect 4638 406 4646 414
rect 4652 406 4660 414
rect 4666 406 4674 414
rect 4972 616 4980 624
rect 4956 596 4964 604
rect 4972 536 4980 544
rect 4956 516 4964 524
rect 4972 496 4980 504
rect 5052 696 5060 704
rect 5068 656 5076 664
rect 5548 1036 5556 1044
rect 5548 1016 5556 1024
rect 5628 1016 5636 1024
rect 5676 1016 5684 1024
rect 5644 956 5652 964
rect 5580 916 5588 924
rect 5628 916 5636 924
rect 5676 916 5684 924
rect 5532 896 5540 904
rect 5628 896 5636 904
rect 5612 876 5620 884
rect 5660 876 5668 884
rect 5548 856 5556 864
rect 5516 796 5524 804
rect 5468 736 5476 744
rect 5532 736 5540 744
rect 5212 696 5220 704
rect 5292 696 5300 704
rect 5436 696 5444 704
rect 5452 696 5460 704
rect 5052 636 5060 644
rect 5100 636 5108 644
rect 5116 636 5124 644
rect 5116 576 5124 584
rect 5164 576 5172 584
rect 5068 556 5076 564
rect 5068 496 5076 504
rect 5020 476 5028 484
rect 5068 456 5076 464
rect 5132 536 5140 544
rect 5260 676 5268 684
rect 5340 676 5348 684
rect 5516 716 5524 724
rect 5500 696 5508 704
rect 5660 696 5668 704
rect 5452 676 5460 684
rect 5548 676 5556 684
rect 5228 656 5236 664
rect 5404 656 5412 664
rect 5324 636 5332 644
rect 5196 616 5204 624
rect 5212 616 5220 624
rect 5212 576 5220 584
rect 5196 536 5204 544
rect 5132 496 5140 504
rect 5180 496 5188 504
rect 5100 456 5108 464
rect 5084 436 5092 444
rect 5148 436 5156 444
rect 5100 416 5108 424
rect 4476 336 4484 344
rect 4908 336 4916 344
rect 4956 336 4964 344
rect 5068 336 5076 344
rect 4572 316 4580 324
rect 4604 316 4612 324
rect 4780 316 4788 324
rect 4620 296 4628 304
rect 4908 296 4916 304
rect 4940 296 4948 304
rect 4876 276 4884 284
rect 4300 256 4308 264
rect 4444 256 4452 264
rect 4524 256 4532 264
rect 4252 236 4260 244
rect 3788 156 3796 164
rect 3868 156 3876 164
rect 4140 156 4148 164
rect 3548 116 3556 124
rect 3660 116 3668 124
rect 3708 96 3716 104
rect 3532 36 3540 44
rect 3564 36 3572 44
rect 3500 16 3508 24
rect 3532 16 3540 24
rect 3788 136 3796 144
rect 3852 136 3860 144
rect 3740 116 3748 124
rect 4044 136 4052 144
rect 3836 116 3844 124
rect 3932 116 3940 124
rect 3788 96 3796 104
rect 4124 36 4132 44
rect 4476 236 4484 244
rect 4316 156 4324 164
rect 4364 156 4372 164
rect 4428 156 4436 164
rect 4252 136 4260 144
rect 4300 136 4308 144
rect 4364 136 4372 144
rect 4380 136 4388 144
rect 4284 96 4292 104
rect 4252 36 4260 44
rect 4460 136 4468 144
rect 4636 236 4644 244
rect 4588 216 4596 224
rect 4812 236 4820 244
rect 4524 136 4532 144
rect 4620 136 4628 144
rect 4780 136 4788 144
rect 4860 196 4868 204
rect 4924 276 4932 284
rect 4876 176 4884 184
rect 4924 176 4932 184
rect 5036 296 5044 304
rect 5132 316 5140 324
rect 5164 316 5172 324
rect 5180 316 5188 324
rect 5004 276 5012 284
rect 5036 276 5044 284
rect 5084 276 5092 284
rect 4988 256 4996 264
rect 4972 236 4980 244
rect 4844 156 4852 164
rect 4892 156 4900 164
rect 4956 156 4964 164
rect 4988 176 4996 184
rect 4748 118 4756 124
rect 4748 116 4756 118
rect 4828 116 4836 124
rect 4892 116 4900 124
rect 5004 116 5012 124
rect 5052 256 5060 264
rect 5340 616 5348 624
rect 5500 596 5508 604
rect 5484 556 5492 564
rect 5532 556 5540 564
rect 5356 536 5364 544
rect 5420 516 5428 524
rect 5388 496 5396 504
rect 5500 516 5508 524
rect 5724 1116 5732 1124
rect 5708 1096 5716 1104
rect 5740 1096 5748 1104
rect 5708 996 5716 1004
rect 5708 956 5716 964
rect 5740 916 5748 924
rect 5708 716 5716 724
rect 5692 576 5700 584
rect 5580 536 5588 544
rect 5580 516 5588 524
rect 5644 516 5652 524
rect 5468 476 5476 484
rect 5516 476 5524 484
rect 5308 436 5316 444
rect 5324 436 5332 444
rect 5244 396 5252 404
rect 5244 356 5252 364
rect 5148 296 5156 304
rect 5228 296 5236 304
rect 5212 276 5220 284
rect 5132 196 5140 204
rect 5356 396 5364 404
rect 5420 396 5428 404
rect 5260 336 5268 344
rect 5340 316 5348 324
rect 5324 296 5332 304
rect 5404 336 5412 344
rect 5388 316 5396 324
rect 5404 316 5412 324
rect 5596 496 5604 504
rect 5628 496 5636 504
rect 5612 476 5620 484
rect 5580 436 5588 444
rect 5564 416 5572 424
rect 5436 356 5444 364
rect 5452 316 5460 324
rect 5516 316 5524 324
rect 5868 1396 5876 1404
rect 5852 1356 5860 1364
rect 6028 2016 6036 2024
rect 6028 1856 6036 1864
rect 6028 1816 6036 1824
rect 6092 2096 6100 2104
rect 6076 2076 6084 2084
rect 6124 2136 6132 2144
rect 6076 2036 6084 2044
rect 6108 2036 6116 2044
rect 6060 1996 6068 2004
rect 6076 1996 6084 2004
rect 6108 1976 6116 1984
rect 6060 1956 6068 1964
rect 6140 2016 6148 2024
rect 6124 1956 6132 1964
rect 6172 2216 6180 2224
rect 6236 2656 6244 2664
rect 6236 2556 6244 2564
rect 6236 2356 6244 2364
rect 6236 2336 6244 2344
rect 6252 2216 6260 2224
rect 6236 2176 6244 2184
rect 6204 2156 6212 2164
rect 6220 2156 6228 2164
rect 6188 2136 6196 2144
rect 6172 2116 6180 2124
rect 6204 2116 6212 2124
rect 6220 2116 6228 2124
rect 6172 2016 6180 2024
rect 6172 1916 6180 1924
rect 6172 1896 6180 1904
rect 6044 1736 6052 1744
rect 6012 1676 6020 1684
rect 6092 1656 6100 1664
rect 6044 1636 6052 1644
rect 6076 1636 6084 1644
rect 5948 1496 5956 1504
rect 5996 1496 6004 1504
rect 6188 1876 6196 1884
rect 6156 1856 6164 1864
rect 6188 1836 6196 1844
rect 6156 1696 6164 1704
rect 6220 2036 6228 2044
rect 6236 1996 6244 2004
rect 6236 1896 6244 1904
rect 6236 1856 6244 1864
rect 6236 1736 6244 1744
rect 6252 1596 6260 1604
rect 6204 1576 6212 1584
rect 6236 1576 6244 1584
rect 6172 1556 6180 1564
rect 5916 1476 5924 1484
rect 6044 1476 6052 1484
rect 6012 1436 6020 1444
rect 5948 1416 5956 1424
rect 5916 1376 5924 1384
rect 5996 1376 6004 1384
rect 6108 1436 6116 1444
rect 5868 1316 5876 1324
rect 5804 1296 5812 1304
rect 5900 1296 5908 1304
rect 5916 1116 5924 1124
rect 5788 1096 5796 1104
rect 5852 1056 5860 1064
rect 5964 1316 5972 1324
rect 6012 1316 6020 1324
rect 6012 1296 6020 1304
rect 6044 1296 6052 1304
rect 6012 1256 6020 1264
rect 5980 1076 5988 1084
rect 6108 1102 6116 1104
rect 6108 1096 6116 1102
rect 6076 1076 6084 1084
rect 6044 1036 6052 1044
rect 6204 1036 6212 1044
rect 6028 976 6036 984
rect 6092 976 6100 984
rect 6156 976 6164 984
rect 5964 936 5972 944
rect 5996 936 6004 944
rect 5852 918 5860 924
rect 5852 916 5860 918
rect 5788 896 5796 904
rect 5772 736 5780 744
rect 5916 776 5924 784
rect 5884 736 5892 744
rect 5916 716 5924 724
rect 5820 696 5828 704
rect 5868 636 5876 644
rect 5804 596 5812 604
rect 5852 596 5860 604
rect 5836 536 5844 544
rect 5692 516 5700 524
rect 5740 516 5748 524
rect 5708 436 5716 444
rect 5676 416 5684 424
rect 5612 396 5620 404
rect 5628 356 5636 364
rect 5612 296 5620 304
rect 5644 336 5652 344
rect 5500 276 5508 284
rect 5532 276 5540 284
rect 5548 276 5556 284
rect 5580 276 5588 284
rect 5436 236 5444 244
rect 5100 176 5108 184
rect 5132 176 5140 184
rect 5308 176 5316 184
rect 5148 156 5156 164
rect 5196 156 5204 164
rect 5260 156 5268 164
rect 5404 216 5412 224
rect 5068 116 5076 124
rect 5228 116 5236 124
rect 5340 116 5348 124
rect 5468 176 5476 184
rect 5548 196 5556 204
rect 5484 156 5492 164
rect 5436 116 5444 124
rect 5468 116 5476 124
rect 4428 96 4436 104
rect 4972 96 4980 104
rect 5084 96 5092 104
rect 5308 96 5316 104
rect 5340 96 5348 104
rect 5420 96 5428 104
rect 5452 96 5460 104
rect 5660 276 5668 284
rect 5660 256 5668 264
rect 5676 256 5684 264
rect 5644 156 5652 164
rect 5676 176 5684 184
rect 5772 476 5780 484
rect 5740 356 5748 364
rect 6188 916 6196 924
rect 5980 896 5988 904
rect 6092 896 6100 904
rect 6140 896 6148 904
rect 6204 876 6212 884
rect 5996 776 6004 784
rect 6188 736 6196 744
rect 6172 696 6180 704
rect 6172 656 6180 664
rect 6236 1016 6244 1024
rect 6236 936 6244 944
rect 6236 716 6244 724
rect 5964 636 5972 644
rect 5948 616 5956 624
rect 5932 576 5940 584
rect 5916 536 5924 544
rect 5820 336 5828 344
rect 5916 336 5924 344
rect 5756 296 5764 304
rect 5820 296 5828 304
rect 5740 216 5748 224
rect 5804 196 5812 204
rect 5612 116 5620 124
rect 5708 116 5716 124
rect 5772 116 5780 124
rect 5564 96 5572 104
rect 5628 96 5636 104
rect 5916 296 5924 304
rect 5900 276 5908 284
rect 5884 256 5892 264
rect 5932 256 5940 264
rect 5916 236 5924 244
rect 5868 196 5876 204
rect 5964 276 5972 284
rect 6172 496 6180 504
rect 6012 336 6020 344
rect 5996 296 6004 304
rect 5996 256 6004 264
rect 6108 256 6116 264
rect 5932 156 5940 164
rect 6220 656 6228 664
rect 6220 636 6228 644
rect 6220 516 6228 524
rect 6204 496 6212 504
rect 6236 456 6244 464
rect 6204 356 6212 364
rect 6124 176 6132 184
rect 5996 136 6004 144
rect 5932 116 5940 124
rect 5964 96 5972 104
rect 6028 96 6036 104
rect 5372 76 5380 84
rect 5548 76 5556 84
rect 5596 76 5604 84
rect 5612 76 5620 84
rect 5820 76 5828 84
rect 4844 16 4852 24
rect 5916 16 5924 24
rect 4638 6 4646 14
rect 4652 6 4660 14
rect 4666 6 4674 14
rect 6156 196 6164 204
rect 6220 316 6228 324
rect 6252 316 6260 324
rect 6156 176 6164 184
rect 6220 156 6228 164
rect 6172 136 6180 144
rect 6172 116 6180 124
rect 6172 16 6180 24
<< metal3 >>
rect 3112 5814 3160 5816
rect 3112 5806 3116 5814
rect 3126 5806 3132 5814
rect 3140 5806 3146 5814
rect 3156 5806 3160 5814
rect 3112 5804 3160 5806
rect 468 5797 492 5803
rect 500 5797 828 5803
rect 1300 5797 1548 5803
rect 3044 5797 3052 5803
rect -19 5777 -13 5783
rect 676 5777 1020 5783
rect 1092 5777 3228 5783
rect 3236 5777 3356 5783
rect 3364 5777 3420 5783
rect 4916 5777 5004 5783
rect 5012 5777 5036 5783
rect 68 5757 124 5763
rect 141 5757 300 5763
rect -19 5737 -13 5743
rect 141 5743 147 5757
rect 660 5757 956 5763
rect 1156 5757 1196 5763
rect 1604 5757 1772 5763
rect 1780 5757 1820 5763
rect 1860 5757 1932 5763
rect 1988 5757 2156 5763
rect 2164 5757 2220 5763
rect 2676 5757 2716 5763
rect 2788 5757 3020 5763
rect 3556 5757 3628 5763
rect 3860 5757 4124 5763
rect 4132 5757 4172 5763
rect 4404 5757 4444 5763
rect 4452 5757 4588 5763
rect 4996 5757 5148 5763
rect 5412 5757 5452 5763
rect 5460 5757 5596 5763
rect 5844 5757 5996 5763
rect 6148 5757 6172 5763
rect 132 5737 147 5743
rect 164 5737 220 5743
rect 228 5737 284 5743
rect 292 5737 364 5743
rect 404 5737 540 5743
rect 804 5737 956 5743
rect 1028 5737 1052 5743
rect 1076 5737 1116 5743
rect 1140 5737 1388 5743
rect 1412 5737 1724 5743
rect 1732 5737 1900 5743
rect 1908 5737 2092 5743
rect 2132 5737 2652 5743
rect 2708 5737 2796 5743
rect 3220 5737 3292 5743
rect 3620 5737 3804 5743
rect 3892 5737 4060 5743
rect 4068 5737 4124 5743
rect 4148 5737 4220 5743
rect 4244 5737 4444 5743
rect 4724 5737 5164 5743
rect 5252 5737 5452 5743
rect 5908 5737 5916 5743
rect 36 5717 76 5723
rect 84 5717 140 5723
rect 212 5717 252 5723
rect 452 5717 508 5723
rect 548 5717 572 5723
rect 788 5717 812 5723
rect 820 5717 908 5723
rect 1012 5717 1468 5723
rect 1476 5717 1628 5723
rect 1652 5717 1916 5723
rect 1940 5717 1996 5723
rect 2052 5717 2140 5723
rect 2148 5717 2204 5723
rect 2221 5717 2300 5723
rect 52 5697 76 5703
rect 372 5697 396 5703
rect 500 5697 540 5703
rect 548 5697 588 5703
rect 852 5697 924 5703
rect 964 5697 1132 5703
rect 1220 5697 1324 5703
rect 1524 5697 1676 5703
rect 1684 5697 1868 5703
rect 1876 5697 2076 5703
rect 2221 5703 2227 5717
rect 2308 5717 2332 5723
rect 2580 5717 2620 5723
rect 2628 5717 2780 5723
rect 3092 5717 3260 5723
rect 3268 5717 3388 5723
rect 3524 5717 3596 5723
rect 3604 5717 3692 5723
rect 4100 5717 4748 5723
rect 4756 5717 4924 5723
rect 5076 5717 5116 5723
rect 5924 5717 5996 5723
rect 2196 5697 2227 5703
rect 2260 5697 2348 5703
rect 2356 5697 2364 5703
rect 2500 5697 2684 5703
rect 2692 5697 2748 5703
rect 2996 5697 3212 5703
rect 3300 5697 3340 5703
rect 3476 5697 3548 5703
rect 4436 5697 4508 5703
rect 4532 5697 4604 5703
rect 4772 5697 4844 5703
rect 4852 5697 4892 5703
rect 4980 5697 5020 5703
rect 5444 5697 5516 5703
rect 5540 5697 5612 5703
rect 5908 5697 6060 5703
rect 6132 5697 6172 5703
rect 612 5677 844 5683
rect 980 5677 1420 5683
rect 1716 5677 1756 5683
rect 1764 5677 1804 5683
rect 1892 5677 1948 5683
rect 1956 5677 2044 5683
rect 2068 5677 2124 5683
rect 2132 5677 2268 5683
rect 2276 5677 2396 5683
rect 2420 5677 2924 5683
rect 2932 5677 3132 5683
rect 3252 5677 3404 5683
rect 4564 5677 4732 5683
rect 4820 5677 5100 5683
rect 6036 5677 6188 5683
rect 324 5657 1084 5663
rect 1108 5657 1372 5663
rect 1780 5657 2284 5663
rect 2292 5657 2380 5663
rect 2628 5657 2812 5663
rect 4276 5657 4956 5663
rect 4964 5657 5052 5663
rect 916 5637 1020 5643
rect 1076 5637 1132 5643
rect 1140 5637 1148 5643
rect 1220 5637 2428 5643
rect 2436 5637 2556 5643
rect 2564 5637 2572 5643
rect 2724 5637 2860 5643
rect 5236 5637 5276 5643
rect 1300 5617 1340 5623
rect 1796 5617 1852 5623
rect 1860 5617 1916 5623
rect 2548 5617 2572 5623
rect 2756 5617 2876 5623
rect 1560 5614 1608 5616
rect 1560 5606 1564 5614
rect 1574 5606 1580 5614
rect 1588 5606 1594 5614
rect 1604 5606 1608 5614
rect 1560 5604 1608 5606
rect 4632 5614 4680 5616
rect 4632 5606 4636 5614
rect 4646 5606 4652 5614
rect 4660 5606 4666 5614
rect 4676 5606 4680 5614
rect 4632 5604 4680 5606
rect 196 5597 236 5603
rect 244 5597 284 5603
rect 1060 5597 1123 5603
rect 212 5577 748 5583
rect 852 5577 1100 5583
rect 1117 5583 1123 5597
rect 1172 5597 1356 5603
rect 1380 5597 1500 5603
rect 3732 5597 4284 5603
rect 1117 5577 1420 5583
rect 1524 5577 1548 5583
rect 1588 5577 1884 5583
rect 2212 5577 2284 5583
rect 2372 5577 2444 5583
rect 3604 5577 3884 5583
rect 4740 5577 4796 5583
rect 5044 5577 5324 5583
rect 5364 5577 5420 5583
rect 5428 5577 5436 5583
rect 5556 5577 5932 5583
rect 52 5557 716 5563
rect 788 5557 3244 5563
rect 3780 5557 3884 5563
rect 3892 5557 5404 5563
rect 5604 5557 5788 5563
rect 5812 5557 5932 5563
rect 100 5537 236 5543
rect 356 5537 460 5543
rect 740 5537 908 5543
rect 996 5537 1340 5543
rect 1364 5537 1436 5543
rect 1444 5537 1980 5543
rect 1988 5537 2044 5543
rect 2148 5537 2332 5543
rect 2340 5537 2380 5543
rect 2804 5537 2860 5543
rect 2884 5537 2908 5543
rect 2916 5537 2972 5543
rect 2980 5537 3004 5543
rect 3236 5537 3260 5543
rect 3348 5537 3436 5543
rect 4228 5537 4252 5543
rect 4260 5537 4300 5543
rect 4308 5537 4380 5543
rect 4612 5537 4892 5543
rect 4900 5537 4940 5543
rect 5140 5537 5196 5543
rect 5204 5537 5228 5543
rect 5300 5537 5356 5543
rect 5389 5537 5452 5543
rect 5389 5524 5395 5537
rect 5492 5537 5548 5543
rect 5556 5537 5692 5543
rect 5988 5537 6076 5543
rect 6244 5537 6252 5543
rect 228 5517 268 5523
rect 1028 5517 1052 5523
rect 1236 5517 1260 5523
rect 1300 5517 1356 5523
rect 1476 5517 1932 5523
rect 2116 5517 2188 5523
rect 2308 5517 2428 5523
rect 2436 5517 2716 5523
rect 2996 5517 3116 5523
rect 3220 5517 3276 5523
rect 3492 5517 3628 5523
rect 3636 5517 3740 5523
rect 4116 5517 4284 5523
rect 4292 5517 4412 5523
rect 4420 5517 4476 5523
rect 4500 5517 4604 5523
rect 4916 5517 5388 5523
rect 5460 5517 5516 5523
rect 5524 5517 5708 5523
rect 196 5497 380 5503
rect 388 5497 428 5503
rect 500 5497 668 5503
rect 884 5497 940 5503
rect 964 5497 988 5503
rect 1284 5497 1388 5503
rect 1412 5497 1580 5503
rect 1620 5497 1772 5503
rect 2180 5497 2284 5503
rect 2372 5497 2396 5503
rect 2404 5497 2636 5503
rect 3188 5497 3292 5503
rect 3300 5497 3356 5503
rect 3412 5497 3452 5503
rect 3684 5497 3708 5503
rect 3876 5497 3932 5503
rect 4052 5497 4156 5503
rect 4324 5497 4716 5503
rect 4756 5497 4908 5503
rect 4916 5497 4956 5503
rect 5044 5497 5068 5503
rect 5108 5497 5212 5503
rect 5332 5497 5372 5503
rect 5380 5497 5468 5503
rect 5684 5497 5836 5503
rect 6100 5497 6156 5503
rect 180 5477 396 5483
rect 404 5477 444 5483
rect 612 5477 716 5483
rect 724 5477 796 5483
rect 1300 5477 1484 5483
rect 1524 5477 1660 5483
rect 1700 5477 1756 5483
rect 2100 5477 2348 5483
rect 2388 5477 2572 5483
rect 2628 5477 2668 5483
rect 2708 5477 2828 5483
rect 2836 5477 2940 5483
rect 2948 5477 3052 5483
rect 3284 5477 3308 5483
rect 3332 5477 3388 5483
rect 3396 5477 3436 5483
rect 3940 5477 3948 5483
rect 3988 5477 4060 5483
rect 4068 5477 4124 5483
rect 4132 5477 4188 5483
rect 4372 5477 4428 5483
rect 5028 5477 5084 5483
rect 5092 5477 5164 5483
rect 5204 5477 5596 5483
rect 5796 5477 6060 5483
rect 6164 5477 6172 5483
rect 260 5457 332 5463
rect 516 5457 620 5463
rect 804 5457 908 5463
rect 1124 5457 1148 5463
rect 1284 5457 1340 5463
rect 1396 5457 1516 5463
rect 1636 5457 1916 5463
rect 1789 5444 1795 5457
rect 1956 5457 2092 5463
rect 2100 5457 2124 5463
rect 2228 5457 2380 5463
rect 2596 5457 2812 5463
rect 3188 5457 3420 5463
rect 3949 5463 3955 5476
rect 3949 5457 3996 5463
rect 4164 5457 4572 5463
rect 4580 5457 4604 5463
rect 4980 5457 5228 5463
rect 5252 5457 5340 5463
rect 5364 5457 5388 5463
rect 5412 5457 5612 5463
rect 5732 5457 5900 5463
rect 5908 5457 6012 5463
rect 148 5437 268 5443
rect 292 5437 380 5443
rect 404 5437 412 5443
rect 468 5437 524 5443
rect 596 5437 1004 5443
rect 1012 5437 1036 5443
rect 1156 5437 1324 5443
rect 1540 5437 1708 5443
rect 1844 5437 1900 5443
rect 1908 5437 1996 5443
rect 2436 5437 2860 5443
rect 2868 5437 2956 5443
rect 2964 5437 3020 5443
rect 3700 5437 3747 5443
rect 244 5417 348 5423
rect 452 5417 540 5423
rect 996 5417 1420 5423
rect 1476 5417 1628 5423
rect 1636 5417 1644 5423
rect 1652 5417 1868 5423
rect 2516 5417 2684 5423
rect 2692 5417 2876 5423
rect 2884 5417 2924 5423
rect 2932 5417 3068 5423
rect 3741 5423 3747 5437
rect 3764 5437 3804 5443
rect 3956 5437 4092 5443
rect 4100 5437 4268 5443
rect 4276 5437 4380 5443
rect 4388 5437 4524 5443
rect 4644 5437 4780 5443
rect 4852 5437 4876 5443
rect 5412 5437 5532 5443
rect 5540 5437 5564 5443
rect 3741 5417 3900 5423
rect 3908 5417 3996 5423
rect 4932 5417 4956 5423
rect 4964 5417 4988 5423
rect 5524 5417 5804 5423
rect 3112 5414 3160 5416
rect 3112 5406 3116 5414
rect 3126 5406 3132 5414
rect 3140 5406 3146 5414
rect 3156 5406 3160 5414
rect 3112 5404 3160 5406
rect -19 5397 -13 5403
rect 180 5397 348 5403
rect 612 5397 828 5403
rect 836 5397 972 5403
rect 1012 5397 1100 5403
rect 1108 5397 1260 5403
rect 2100 5397 2748 5403
rect 5652 5397 5900 5403
rect 20 5377 28 5383
rect 36 5377 444 5383
rect 468 5377 652 5383
rect 852 5377 1132 5383
rect 1252 5377 1260 5383
rect 2324 5377 2476 5383
rect 2484 5377 2540 5383
rect 2580 5377 2812 5383
rect 2836 5377 3180 5383
rect 3220 5377 3372 5383
rect 3572 5377 3580 5383
rect 3604 5377 3932 5383
rect 4068 5377 4316 5383
rect 4916 5377 4972 5383
rect 5620 5377 5660 5383
rect 6116 5377 6172 5383
rect -19 5357 -13 5363
rect 148 5357 220 5363
rect 237 5357 492 5363
rect 20 5337 28 5343
rect 237 5343 243 5357
rect 724 5357 1068 5363
rect 1140 5357 1196 5363
rect 1204 5357 1612 5363
rect 1700 5357 1724 5363
rect 2276 5357 2284 5363
rect 2372 5357 2412 5363
rect 2628 5357 2716 5363
rect 2804 5357 2844 5363
rect 2852 5357 2892 5363
rect 2900 5357 2956 5363
rect 3108 5357 3340 5363
rect 3748 5357 4092 5363
rect 4100 5357 4140 5363
rect 4212 5357 4284 5363
rect 4900 5357 4924 5363
rect 5860 5357 5948 5363
rect 5997 5363 6003 5376
rect 5988 5357 6003 5363
rect 6068 5357 6220 5363
rect 36 5337 243 5343
rect 260 5337 284 5343
rect 436 5337 492 5343
rect 500 5337 540 5343
rect 740 5337 844 5343
rect 916 5337 1212 5343
rect 1220 5337 1308 5343
rect 1428 5337 1532 5343
rect 1652 5337 1692 5343
rect 2052 5337 2332 5343
rect 2340 5337 2396 5343
rect 2516 5337 3020 5343
rect 3028 5337 3100 5343
rect 3204 5337 3228 5343
rect 3268 5337 3324 5343
rect 3508 5337 3516 5343
rect 3796 5337 3884 5343
rect 3892 5337 3980 5343
rect 4308 5337 4460 5343
rect 4596 5337 4732 5343
rect 4900 5337 5228 5343
rect 5236 5337 5292 5343
rect 5348 5337 5420 5343
rect 5428 5337 5532 5343
rect 5556 5337 5692 5343
rect 5700 5337 5788 5343
rect 5844 5337 6012 5343
rect -19 5317 -13 5323
rect 52 5317 156 5323
rect 308 5317 412 5323
rect 452 5317 556 5323
rect 628 5317 828 5323
rect 900 5317 1036 5323
rect 1044 5317 1068 5323
rect 1124 5317 1180 5323
rect 1316 5317 1356 5323
rect 1428 5317 1468 5323
rect 1700 5317 1820 5323
rect 1828 5317 1868 5323
rect 1876 5317 1916 5323
rect 2148 5317 2204 5323
rect 2212 5317 2268 5323
rect 2372 5317 2556 5323
rect 2564 5317 2764 5323
rect 3012 5317 3068 5323
rect 3076 5317 3308 5323
rect 3316 5317 3356 5323
rect 3428 5317 3628 5323
rect 3700 5317 3740 5323
rect 3780 5317 3820 5323
rect 3853 5317 4124 5323
rect 84 5297 252 5303
rect 404 5297 444 5303
rect 484 5297 508 5303
rect 516 5297 572 5303
rect 1092 5297 1164 5303
rect 1204 5297 1340 5303
rect 1348 5297 1452 5303
rect 1492 5297 1596 5303
rect 1828 5297 1900 5303
rect 1908 5297 1948 5303
rect 1988 5297 2108 5303
rect 2180 5297 2316 5303
rect 2324 5297 2380 5303
rect 2660 5297 2700 5303
rect 2708 5297 2780 5303
rect 2804 5297 2860 5303
rect 2868 5297 2908 5303
rect 2916 5297 2940 5303
rect 3060 5297 3180 5303
rect 3284 5297 3404 5303
rect 3853 5303 3859 5317
rect 4132 5317 4188 5323
rect 4228 5317 4316 5323
rect 4484 5317 4508 5323
rect 4580 5317 4684 5323
rect 4804 5317 4908 5323
rect 4980 5317 5036 5323
rect 5076 5317 5116 5323
rect 5124 5317 5164 5323
rect 5236 5317 5308 5323
rect 5476 5317 5612 5323
rect 5716 5317 5756 5323
rect 5828 5317 5884 5323
rect 5924 5317 5932 5323
rect 6020 5317 6044 5323
rect 6132 5317 6188 5323
rect 3492 5297 3859 5303
rect 3876 5297 4108 5303
rect 4116 5297 4156 5303
rect 4292 5297 4556 5303
rect 4564 5297 4700 5303
rect 4868 5297 4892 5303
rect 4964 5297 5100 5303
rect 5108 5297 5132 5303
rect 5140 5297 5180 5303
rect 5364 5297 5484 5303
rect 5492 5297 5548 5303
rect 5556 5297 5580 5303
rect 5684 5297 5852 5303
rect 6228 5297 6291 5303
rect 628 5277 636 5283
rect 1076 5277 1292 5283
rect 1380 5277 1404 5283
rect 1412 5277 1500 5283
rect 1524 5277 1740 5283
rect 1780 5277 1804 5283
rect 1812 5277 1852 5283
rect 2036 5277 2076 5283
rect 2164 5277 2188 5283
rect 2196 5277 2284 5283
rect 2500 5277 2668 5283
rect 2676 5277 2700 5283
rect 2724 5277 2764 5283
rect 2772 5277 2796 5283
rect 2916 5277 2972 5283
rect 3300 5277 3324 5283
rect 3508 5277 3692 5283
rect 3700 5277 3836 5283
rect 5172 5277 5244 5283
rect 5476 5277 5532 5283
rect 5668 5277 5740 5283
rect 5812 5277 5852 5283
rect 1060 5257 1356 5263
rect 1364 5257 1436 5263
rect 1444 5257 1564 5263
rect 1572 5257 1708 5263
rect 1716 5257 1756 5263
rect 2020 5257 2092 5263
rect 2100 5257 2172 5263
rect 4724 5257 4956 5263
rect 5092 5257 5132 5263
rect 5140 5257 5212 5263
rect 5444 5257 5500 5263
rect 5508 5257 5612 5263
rect 5748 5257 5772 5263
rect 36 5237 60 5243
rect 244 5237 396 5243
rect 1444 5237 1964 5243
rect 1972 5237 1996 5243
rect 2004 5237 2236 5243
rect 2244 5237 2252 5243
rect 3812 5237 3852 5243
rect 3860 5237 4044 5243
rect 4468 5237 5340 5243
rect 5572 5237 5628 5243
rect 6196 5237 6252 5243
rect 6285 5237 6291 5243
rect 1700 5217 1724 5223
rect 4932 5217 5020 5223
rect 5028 5217 5180 5223
rect 5588 5217 6188 5223
rect 1560 5214 1608 5216
rect 1560 5206 1564 5214
rect 1574 5206 1580 5214
rect 1588 5206 1594 5214
rect 1604 5206 1608 5214
rect 1560 5204 1608 5206
rect 4632 5214 4680 5216
rect 4632 5206 4636 5214
rect 4646 5206 4652 5214
rect 4660 5206 4666 5214
rect 4676 5206 4680 5214
rect 4632 5204 4680 5206
rect 3924 5197 3948 5203
rect 5156 5197 5452 5203
rect 5460 5197 5516 5203
rect 836 5177 1996 5183
rect 3428 5177 3564 5183
rect 3924 5177 3948 5183
rect 4276 5177 4492 5183
rect 4500 5177 4524 5183
rect 4996 5177 5436 5183
rect 5444 5177 5484 5183
rect 3540 5157 3612 5163
rect 3748 5157 4188 5163
rect 4372 5157 4396 5163
rect 4484 5157 4908 5163
rect 4916 5157 4940 5163
rect 4948 5157 5020 5163
rect 5252 5157 5676 5163
rect 5684 5157 5740 5163
rect 836 5137 892 5143
rect 1076 5137 1180 5143
rect 1780 5137 2140 5143
rect 3060 5137 3148 5143
rect 3156 5137 3244 5143
rect 3444 5137 3484 5143
rect 3492 5137 3532 5143
rect 3556 5137 3708 5143
rect 3876 5137 3932 5143
rect 4308 5137 4700 5143
rect 4708 5137 4748 5143
rect 4756 5137 4828 5143
rect 5364 5137 5500 5143
rect 5508 5137 5548 5143
rect 5748 5137 6204 5143
rect 276 5117 380 5123
rect 596 5117 716 5123
rect 772 5117 956 5123
rect 1044 5117 1244 5123
rect 1332 5117 1468 5123
rect 1476 5117 1740 5123
rect 1924 5117 1948 5123
rect 3268 5117 3324 5123
rect 3380 5117 3404 5123
rect 3460 5117 3468 5123
rect 3476 5117 3644 5123
rect 3652 5117 3708 5123
rect 3796 5117 3884 5123
rect 4084 5117 4140 5123
rect 4212 5117 4300 5123
rect 4340 5117 4428 5123
rect 4436 5117 4460 5123
rect 4548 5117 4716 5123
rect 4724 5117 4764 5123
rect 4772 5117 4812 5123
rect 5220 5117 5244 5123
rect 5284 5117 5420 5123
rect 5428 5117 5516 5123
rect 5620 5117 5708 5123
rect 5828 5117 5868 5123
rect 5956 5117 5964 5123
rect 228 5097 284 5103
rect 292 5097 332 5103
rect 436 5097 476 5103
rect 708 5097 828 5103
rect 868 5097 956 5103
rect 973 5097 1004 5103
rect 84 5077 268 5083
rect 452 5077 492 5083
rect 756 5077 908 5083
rect 973 5083 979 5097
rect 1108 5097 1372 5103
rect 1428 5097 1628 5103
rect 1636 5097 1676 5103
rect 1828 5097 1916 5103
rect 1972 5097 1996 5103
rect 2004 5097 2060 5103
rect 2068 5097 2204 5103
rect 2372 5097 2444 5103
rect 2836 5097 2892 5103
rect 2996 5097 3036 5103
rect 3268 5097 3516 5103
rect 3524 5097 3580 5103
rect 3588 5097 3628 5103
rect 3645 5097 3692 5103
rect 3645 5084 3651 5097
rect 3700 5097 3740 5103
rect 3972 5097 4060 5103
rect 4164 5097 4236 5103
rect 4308 5097 4364 5103
rect 4484 5097 4540 5103
rect 4548 5097 4604 5103
rect 4644 5097 4892 5103
rect 4900 5097 4956 5103
rect 4964 5097 5004 5103
rect 5204 5097 5212 5103
rect 5540 5097 5660 5103
rect 5668 5097 5724 5103
rect 5908 5097 5948 5103
rect 6228 5097 6252 5103
rect 932 5077 979 5083
rect 996 5077 1068 5083
rect 1300 5077 1420 5083
rect 1588 5077 1724 5083
rect 1828 5077 1868 5083
rect 2068 5077 2188 5083
rect 2196 5077 2236 5083
rect 2276 5077 2428 5083
rect 2580 5077 2668 5083
rect 2740 5077 2956 5083
rect 2964 5077 3020 5083
rect 3092 5077 3164 5083
rect 3348 5077 3500 5083
rect 3508 5077 3564 5083
rect 3668 5077 3724 5083
rect 3828 5077 3980 5083
rect 4052 5077 4172 5083
rect 4180 5077 4220 5083
rect 4292 5077 4348 5083
rect 4388 5077 4572 5083
rect 4868 5077 4940 5083
rect 4948 5077 5068 5083
rect 5556 5077 5580 5083
rect 5812 5077 5836 5083
rect 6285 5083 6291 5103
rect 6196 5077 6291 5083
rect 20 5057 76 5063
rect 84 5057 92 5063
rect 324 5057 364 5063
rect 372 5057 444 5063
rect 740 5057 780 5063
rect 900 5057 940 5063
rect 1012 5057 1052 5063
rect 1060 5057 1180 5063
rect 1188 5057 1356 5063
rect 1428 5057 1644 5063
rect 1732 5057 1836 5063
rect 1844 5057 1852 5063
rect 2052 5057 2092 5063
rect 2180 5057 2572 5063
rect 2628 5057 2636 5063
rect 2644 5057 2652 5063
rect 2708 5057 2764 5063
rect 2772 5057 2908 5063
rect 2916 5057 2988 5063
rect 3332 5057 3372 5063
rect 3396 5057 3420 5063
rect 3428 5057 3660 5063
rect 3684 5057 3788 5063
rect 3892 5057 3900 5063
rect 4212 5057 4252 5063
rect 4260 5057 4284 5063
rect 4404 5057 4428 5063
rect 4436 5057 4556 5063
rect 4564 5057 4604 5063
rect 4852 5057 4988 5063
rect 4996 5057 5036 5063
rect 5204 5057 5340 5063
rect -19 5037 -13 5043
rect 196 5037 252 5043
rect 260 5037 380 5043
rect 1060 5037 1100 5043
rect 1172 5037 1308 5043
rect 1716 5037 2316 5043
rect 2324 5037 2412 5043
rect 2436 5037 2588 5043
rect 2596 5037 2684 5043
rect 3572 5037 3772 5043
rect 3780 5037 3852 5043
rect 3892 5037 3964 5043
rect 3988 5037 4236 5043
rect 4356 5037 4572 5043
rect 4740 5037 4796 5043
rect 4804 5037 4876 5043
rect 4884 5037 4988 5043
rect 5044 5037 5084 5043
rect 5140 5037 5228 5043
rect 5236 5037 5260 5043
rect 5300 5037 5340 5043
rect 5780 5037 6076 5043
rect 948 5017 1132 5023
rect 1252 5017 1420 5023
rect 1604 5017 2140 5023
rect 2196 5017 2220 5023
rect 2228 5017 2252 5023
rect 2516 5017 2524 5023
rect 3300 5017 3356 5023
rect 3364 5017 3532 5023
rect 3860 5017 3996 5023
rect 4004 5017 4220 5023
rect 5268 5017 6236 5023
rect 3112 5014 3160 5016
rect 3112 5006 3116 5014
rect 3126 5006 3132 5014
rect 3140 5006 3146 5014
rect 3156 5006 3160 5014
rect 3112 5004 3160 5006
rect 1092 4997 1164 5003
rect 1220 4997 1244 5003
rect 1268 4997 1276 5003
rect 1380 4997 1676 5003
rect 1796 4997 1804 5003
rect 1924 4997 2060 5003
rect 2420 4997 2476 5003
rect 2484 4997 2604 5003
rect 2964 4997 3052 5003
rect 3188 4997 3372 5003
rect 3380 4997 6108 5003
rect 564 4977 924 4983
rect 932 4977 1228 4983
rect 1876 4977 1932 4983
rect 2292 4977 2332 4983
rect 2516 4977 2556 4983
rect 2868 4977 2924 4983
rect 2932 4977 2988 4983
rect 3124 4977 3212 4983
rect 3812 4977 4076 4983
rect 4564 4977 4620 4983
rect 4724 4977 4956 4983
rect 5972 4977 5980 4983
rect 6004 4977 6124 4983
rect 6228 4977 6252 4983
rect 84 4957 220 4963
rect 740 4957 956 4963
rect 1076 4957 1196 4963
rect 1252 4957 1372 4963
rect 1844 4957 1900 4963
rect 1917 4957 1980 4963
rect 116 4937 364 4943
rect 372 4937 412 4943
rect 500 4937 524 4943
rect 980 4937 988 4943
rect 1044 4937 1100 4943
rect 1156 4937 1260 4943
rect 1364 4937 1404 4943
rect 1412 4937 1516 4943
rect 1917 4943 1923 4957
rect 2244 4957 2300 4963
rect 2324 4957 2380 4963
rect 2468 4957 2524 4963
rect 2628 4957 2668 4963
rect 2740 4957 3004 4963
rect 3828 4957 3868 4963
rect 3876 4957 3916 4963
rect 4004 4957 4092 4963
rect 4148 4957 4268 4963
rect 4308 4957 4364 4963
rect 4372 4957 4428 4963
rect 4548 4957 4572 4963
rect 4788 4957 4860 4963
rect 4868 4957 4924 4963
rect 5332 4957 5356 4963
rect 5588 4957 5740 4963
rect 5748 4957 5788 4963
rect 5940 4957 5964 4963
rect 5972 4957 6028 4963
rect 1892 4937 1923 4943
rect 1940 4937 1964 4943
rect 2148 4937 2236 4943
rect 2308 4937 2348 4943
rect 2388 4937 2572 4943
rect 2580 4937 2636 4943
rect 2804 4937 2940 4943
rect 3060 4937 3084 4943
rect 3092 4937 3276 4943
rect 3412 4937 3452 4943
rect 3860 4937 3980 4943
rect 4068 4937 4332 4943
rect 4340 4937 4412 4943
rect 4548 4937 4636 4943
rect 4660 4937 4908 4943
rect 4948 4937 5100 4943
rect 5428 4937 5500 4943
rect 5508 4937 5548 4943
rect 5556 4937 5580 4943
rect 6180 4937 6252 4943
rect 164 4917 204 4923
rect 212 4917 316 4923
rect 676 4917 764 4923
rect 900 4917 1036 4923
rect 1156 4917 1212 4923
rect 1220 4917 1324 4923
rect 1357 4917 1820 4923
rect 132 4897 172 4903
rect 292 4897 332 4903
rect 340 4897 380 4903
rect 516 4897 556 4903
rect 564 4897 700 4903
rect 948 4897 1020 4903
rect 1028 4897 1068 4903
rect 1357 4903 1363 4917
rect 1860 4917 2156 4923
rect 2164 4917 2252 4923
rect 2260 4917 2508 4923
rect 2564 4917 2588 4923
rect 2596 4917 2652 4923
rect 2916 4917 2972 4923
rect 3412 4917 3468 4923
rect 3540 4917 3580 4923
rect 3796 4917 3836 4923
rect 3908 4917 3948 4923
rect 3956 4917 4028 4923
rect 4052 4917 4092 4923
rect 4148 4917 4204 4923
rect 4260 4917 4316 4923
rect 4324 4917 4396 4923
rect 4461 4923 4467 4936
rect 4461 4917 4732 4923
rect 4740 4917 4812 4923
rect 5028 4917 5052 4923
rect 5220 4917 5244 4923
rect 5268 4917 5292 4923
rect 5396 4917 5436 4923
rect 5693 4917 5804 4923
rect 5693 4904 5699 4917
rect 5844 4917 5900 4923
rect 5908 4917 5932 4923
rect 6029 4923 6035 4936
rect 5972 4917 6035 4923
rect 1092 4897 1363 4903
rect 1508 4897 1548 4903
rect 2116 4897 2444 4903
rect 2452 4897 2524 4903
rect 2580 4897 2620 4903
rect 2852 4897 2940 4903
rect 2980 4897 3036 4903
rect 3380 4897 3388 4903
rect 3444 4897 3516 4903
rect 3540 4897 3612 4903
rect 3620 4897 3644 4903
rect 3972 4897 4044 4903
rect 4452 4897 4700 4903
rect 4708 4897 4780 4903
rect 4916 4897 4972 4903
rect 4996 4897 5036 4903
rect 5092 4897 5148 4903
rect 5284 4897 5372 4903
rect 5700 4897 5740 4903
rect 5892 4897 5932 4903
rect 5972 4897 6188 4903
rect 6260 4897 6291 4903
rect 1044 4877 1164 4883
rect 1172 4877 1308 4883
rect 1492 4877 1628 4883
rect 2036 4877 2124 4883
rect 2132 4877 2204 4883
rect 2308 4877 2428 4883
rect 2436 4877 2492 4883
rect 2500 4877 2700 4883
rect 2724 4877 2876 4883
rect 3236 4877 3404 4883
rect 3540 4877 3548 4883
rect 3604 4877 3644 4883
rect 3652 4877 3708 4883
rect 4420 4877 4476 4883
rect 4500 4877 4524 4883
rect 4612 4877 4876 4883
rect 5140 4877 5148 4883
rect 5348 4877 5468 4883
rect 5828 4877 5852 4883
rect 5860 4877 5916 4883
rect 6036 4877 6204 4883
rect 6228 4877 6252 4883
rect 756 4857 2044 4863
rect 2820 4857 3180 4863
rect 3188 4857 3212 4863
rect 3236 4857 3500 4863
rect 3508 4857 3676 4863
rect 3684 4857 3740 4863
rect 5044 4857 5404 4863
rect 5412 4857 5452 4863
rect 5956 4857 5996 4863
rect 564 4837 1724 4843
rect 1940 4837 2364 4843
rect 3044 4837 3388 4843
rect 3396 4837 3420 4843
rect 3476 4837 3660 4843
rect 3668 4837 3724 4843
rect 4580 4837 5436 4843
rect 5876 4837 6044 4843
rect 6068 4837 6140 4843
rect 6148 4837 6188 4843
rect 724 4817 780 4823
rect 1380 4817 1452 4823
rect 1988 4817 2140 4823
rect 3508 4817 3772 4823
rect 3780 4817 3852 4823
rect 5444 4817 5596 4823
rect 5780 4817 6220 4823
rect 6285 4817 6291 4823
rect 1560 4814 1608 4816
rect 1560 4806 1564 4814
rect 1574 4806 1580 4814
rect 1588 4806 1594 4814
rect 1604 4806 1608 4814
rect 1560 4804 1608 4806
rect 4632 4814 4680 4816
rect 4632 4806 4636 4814
rect 4646 4806 4652 4814
rect 4660 4806 4666 4814
rect 4676 4806 4680 4814
rect 4632 4804 4680 4806
rect -19 4797 -13 4803
rect 84 4797 124 4803
rect 1124 4797 1196 4803
rect 1332 4797 1484 4803
rect 1988 4797 2124 4803
rect 3380 4797 3404 4803
rect 4836 4797 4988 4803
rect 5204 4797 5292 4803
rect 5988 4797 6060 4803
rect 1412 4777 2076 4783
rect 2532 4777 2700 4783
rect 3652 4777 3788 4783
rect 3796 4777 3884 4783
rect 3892 4777 4012 4783
rect 4324 4777 4796 4783
rect 4804 4777 4844 4783
rect 4852 4777 5020 4783
rect 5748 4777 5891 4783
rect 820 4757 972 4763
rect 1300 4757 1388 4763
rect 1540 4757 1612 4763
rect 1796 4757 2380 4763
rect 2436 4757 2572 4763
rect 2660 4757 2860 4763
rect 3028 4757 3052 4763
rect 3780 4757 4076 4763
rect 4260 4757 4300 4763
rect 4308 4757 4364 4763
rect 4388 4757 4572 4763
rect 4580 4757 4604 4763
rect 5012 4757 5772 4763
rect 5812 4757 5852 4763
rect 5885 4763 5891 4777
rect 5908 4777 5932 4783
rect 5885 4757 5932 4763
rect 5940 4757 6060 4763
rect 948 4737 1324 4743
rect 1332 4737 1388 4743
rect 1460 4737 1660 4743
rect 1668 4737 1756 4743
rect 1780 4737 1836 4743
rect 1844 4737 1884 4743
rect 1908 4737 1996 4743
rect 2468 4737 2508 4743
rect 2596 4737 2620 4743
rect 2852 4737 2908 4743
rect 2964 4737 3052 4743
rect 3364 4737 3500 4743
rect 3508 4737 3564 4743
rect 3764 4737 3836 4743
rect 4068 4737 4316 4743
rect 4324 4737 4380 4743
rect 4484 4737 4556 4743
rect 4564 4737 4620 4743
rect 4996 4737 5116 4743
rect 5252 4737 5516 4743
rect 5524 4737 5644 4743
rect 5764 4737 5820 4743
rect 5828 4737 5836 4743
rect 5940 4737 6156 4743
rect 644 4717 684 4723
rect 900 4717 972 4723
rect 1444 4717 1516 4723
rect 1629 4717 2083 4723
rect 196 4697 332 4703
rect 484 4697 668 4703
rect 948 4697 972 4703
rect 980 4697 1052 4703
rect 1316 4697 1372 4703
rect 1380 4697 1420 4703
rect 1629 4703 1635 4717
rect 1492 4697 1635 4703
rect 1652 4697 1852 4703
rect 1860 4697 1900 4703
rect 1972 4697 2028 4703
rect 2077 4703 2083 4717
rect 2100 4717 2156 4723
rect 2164 4717 2252 4723
rect 2484 4717 2556 4723
rect 2580 4717 2652 4723
rect 2772 4717 2988 4723
rect 3268 4717 3292 4723
rect 3348 4717 3420 4723
rect 3780 4717 3820 4723
rect 3860 4717 3884 4723
rect 3892 4717 4012 4723
rect 4020 4717 4044 4723
rect 4148 4717 4204 4723
rect 4317 4717 4412 4723
rect 2077 4697 2220 4703
rect 2468 4697 2492 4703
rect 2500 4697 2524 4703
rect 2612 4697 2716 4703
rect 2804 4697 2940 4703
rect 2948 4697 3084 4703
rect 3252 4697 3308 4703
rect 3412 4697 3436 4703
rect 3732 4697 3756 4703
rect 3796 4697 3836 4703
rect 3860 4697 3948 4703
rect 4020 4697 4060 4703
rect 4068 4697 4108 4703
rect 4317 4703 4323 4717
rect 4420 4717 4492 4723
rect 4644 4717 5244 4723
rect 5252 4717 5308 4723
rect 5492 4717 5532 4723
rect 5540 4717 5660 4723
rect 5796 4717 5948 4723
rect 5956 4717 6044 4723
rect 6084 4717 6108 4723
rect 4132 4697 4323 4703
rect 4340 4697 4460 4703
rect 4468 4697 4508 4703
rect 4756 4697 4780 4703
rect 5044 4697 5068 4703
rect 5428 4697 5468 4703
rect 5508 4697 5708 4703
rect 5716 4697 5772 4703
rect 5876 4697 5980 4703
rect 6100 4697 6108 4703
rect 6125 4697 6140 4703
rect 6125 4684 6131 4697
rect 6212 4697 6220 4703
rect 164 4677 236 4683
rect 452 4677 652 4683
rect 852 4677 1084 4683
rect 1092 4677 1164 4683
rect 1284 4677 1452 4683
rect 1460 4677 1532 4683
rect 1924 4677 1980 4683
rect 1988 4677 2028 4683
rect 2148 4677 2172 4683
rect 2548 4677 2668 4683
rect 2964 4677 3100 4683
rect 3236 4677 3260 4683
rect 3332 4677 3484 4683
rect 3492 4677 3548 4683
rect 3748 4677 3932 4683
rect 4212 4677 4236 4683
rect 4388 4677 4412 4683
rect 4420 4677 4476 4683
rect 4532 4677 4812 4683
rect 4820 4677 4860 4683
rect 4884 4677 5228 4683
rect 5236 4677 5292 4683
rect 5364 4677 5564 4683
rect 5588 4677 5692 4683
rect 5700 4677 5756 4683
rect 5892 4677 6028 4683
rect 6100 4677 6124 4683
rect 6141 4677 6172 4683
rect 20 4657 108 4663
rect 452 4657 476 4663
rect 516 4657 556 4663
rect 564 4657 668 4663
rect 916 4657 1020 4663
rect 1140 4657 1164 4663
rect 1188 4657 1676 4663
rect 1684 4657 1772 4663
rect 1876 4657 1932 4663
rect 2212 4657 2348 4663
rect 2356 4657 2428 4663
rect 2804 4657 2828 4663
rect 2836 4657 3020 4663
rect 3028 4657 3052 4663
rect 3412 4657 3452 4663
rect 3460 4657 3548 4663
rect 3668 4657 3724 4663
rect 3732 4657 3756 4663
rect 3780 4657 3820 4663
rect 3844 4657 4268 4663
rect 4276 4657 4412 4663
rect 4436 4657 4460 4663
rect 4660 4657 4764 4663
rect 4772 4657 4828 4663
rect 4980 4657 5052 4663
rect 5300 4657 5324 4663
rect 5364 4657 5388 4663
rect 5492 4657 5580 4663
rect 5700 4657 5724 4663
rect 5732 4657 5740 4663
rect 5908 4657 6012 4663
rect 6141 4663 6147 4677
rect 6036 4657 6147 4663
rect 84 4637 140 4643
rect 212 4637 268 4643
rect 500 4637 524 4643
rect 532 4637 652 4643
rect 788 4637 940 4643
rect 1028 4637 1196 4643
rect 1236 4637 1292 4643
rect 1636 4637 1660 4643
rect 2148 4637 2364 4643
rect 2372 4637 2444 4643
rect 3220 4637 3276 4643
rect 3284 4637 3436 4643
rect 3908 4637 4252 4643
rect 4260 4637 4396 4643
rect 4772 4637 4924 4643
rect 4932 4637 5052 4643
rect 5124 4637 5436 4643
rect 5524 4637 5884 4643
rect 276 4617 348 4623
rect 628 4617 876 4623
rect 1172 4617 1292 4623
rect 1476 4617 1516 4623
rect 1524 4617 1644 4623
rect 1652 4617 1804 4623
rect 2468 4617 2659 4623
rect 116 4597 220 4603
rect 836 4597 892 4603
rect 1108 4597 1340 4603
rect 1348 4597 1404 4603
rect 1444 4597 1500 4603
rect 2653 4603 2659 4617
rect 2676 4617 2700 4623
rect 3412 4617 3644 4623
rect 3652 4617 3676 4623
rect 3892 4617 3932 4623
rect 4116 4617 4444 4623
rect 4916 4617 4972 4623
rect 5028 4617 5212 4623
rect 5220 4617 5356 4623
rect 5604 4617 5676 4623
rect 5716 4617 5964 4623
rect 6052 4617 6236 4623
rect 3112 4614 3160 4616
rect 3112 4606 3116 4614
rect 3126 4606 3132 4614
rect 3140 4606 3146 4614
rect 3156 4606 3160 4614
rect 3112 4604 3160 4606
rect 2653 4597 2828 4603
rect 2836 4597 2876 4603
rect 3572 4597 3628 4603
rect 3636 4597 3692 4603
rect 4052 4597 4284 4603
rect 4404 4597 4540 4603
rect 4548 4597 4604 4603
rect 4996 4597 5100 4603
rect 5796 4597 5852 4603
rect 5908 4597 6092 4603
rect -19 4577 12 4583
rect 356 4577 492 4583
rect 500 4577 860 4583
rect 868 4577 972 4583
rect 1332 4577 1596 4583
rect 1604 4577 1724 4583
rect 1748 4577 2188 4583
rect 2196 4577 2284 4583
rect 2397 4577 2620 4583
rect 2397 4564 2403 4577
rect 3188 4577 3228 4583
rect 3268 4577 3612 4583
rect 3764 4577 3852 4583
rect 4068 4577 4140 4583
rect 4244 4577 4492 4583
rect 4596 4577 4924 4583
rect 5092 4577 5116 4583
rect 5124 4577 5164 4583
rect 5492 4577 5980 4583
rect 132 4557 188 4563
rect 580 4557 636 4563
rect 996 4557 1100 4563
rect 1172 4557 1228 4563
rect 1268 4557 1324 4563
rect 1748 4557 1852 4563
rect 1956 4557 2172 4563
rect 2180 4557 2268 4563
rect 2340 4557 2396 4563
rect 2420 4557 2492 4563
rect 2500 4557 2588 4563
rect 2596 4557 2668 4563
rect 3764 4557 3868 4563
rect 4020 4557 4092 4563
rect 4164 4557 4300 4563
rect 4868 4557 5004 4563
rect 5380 4557 5564 4563
rect 5572 4557 5676 4563
rect 5844 4557 6092 4563
rect 6100 4557 6140 4563
rect -19 4537 -13 4543
rect 20 4537 236 4543
rect 468 4537 748 4543
rect 772 4537 876 4543
rect 1428 4537 1628 4543
rect 1636 4537 1932 4543
rect 1940 4537 1996 4543
rect 2068 4537 2108 4543
rect 2324 4537 2412 4543
rect 2788 4537 2924 4543
rect 2932 4537 2972 4543
rect 3076 4537 3276 4543
rect 3652 4537 3884 4543
rect 3940 4537 3980 4543
rect 4100 4537 4124 4543
rect 4132 4537 4188 4543
rect 4196 4537 4252 4543
rect 4292 4537 4316 4543
rect 4404 4537 4476 4543
rect 4724 4537 4828 4543
rect 4836 4537 4908 4543
rect 4916 4537 5020 4543
rect 5149 4537 5228 4543
rect 292 4517 412 4523
rect 484 4517 492 4523
rect 500 4517 716 4523
rect 1236 4517 1916 4523
rect 1924 4517 1980 4523
rect 2036 4517 2076 4523
rect 2084 4517 2124 4523
rect 2276 4517 2540 4523
rect 2548 4517 2572 4523
rect 2580 4517 2652 4523
rect 2820 4517 2860 4523
rect 3060 4517 3324 4523
rect 3476 4517 3500 4523
rect 3588 4517 3612 4523
rect 4548 4517 4572 4523
rect 4724 4517 4796 4523
rect 4804 4517 4876 4523
rect 5149 4523 5155 4537
rect 5252 4537 5308 4543
rect 5412 4537 5452 4543
rect 5620 4537 5724 4543
rect 5732 4537 5756 4543
rect 5844 4537 5868 4543
rect 5972 4537 5996 4543
rect 6068 4537 6124 4543
rect 6164 4537 6204 4543
rect 5140 4517 5155 4523
rect 5236 4517 5260 4523
rect 5300 4517 5372 4523
rect 5572 4517 5644 4523
rect 5876 4517 5916 4523
rect 6084 4517 6108 4523
rect 452 4497 476 4503
rect 564 4497 604 4503
rect 660 4497 684 4503
rect 708 4497 764 4503
rect 948 4497 1036 4503
rect 1044 4497 1052 4503
rect 1348 4497 1420 4503
rect 1476 4497 1500 4503
rect 1764 4497 1836 4503
rect 1844 4497 1900 4503
rect 2084 4497 2476 4503
rect 2484 4497 2524 4503
rect 2532 4497 2556 4503
rect 2788 4497 2812 4503
rect 2948 4497 2988 4503
rect 3060 4497 3084 4503
rect 3172 4497 3244 4503
rect 3252 4497 3372 4503
rect 3380 4497 3388 4503
rect 3428 4497 3452 4503
rect 3812 4497 3948 4503
rect 4148 4497 4220 4503
rect 4596 4497 4620 4503
rect 4708 4497 4764 4503
rect 4868 4497 4908 4503
rect 5108 4497 5276 4503
rect 5396 4497 5596 4503
rect 5732 4497 5900 4503
rect 6100 4497 6124 4503
rect 52 4477 460 4483
rect 548 4477 588 4483
rect 660 4477 684 4483
rect 708 4477 988 4483
rect 996 4477 1084 4483
rect 1316 4477 1740 4483
rect 1812 4477 2060 4483
rect 2100 4477 2156 4483
rect 2164 4477 2476 4483
rect 2660 4477 2732 4483
rect 2740 4477 2908 4483
rect 3028 4477 3052 4483
rect 3060 4477 3148 4483
rect 3284 4477 3308 4483
rect 3348 4477 3516 4483
rect 3524 4477 3532 4483
rect 3540 4477 3628 4483
rect 3956 4477 4172 4483
rect 4180 4477 4236 4483
rect 4772 4477 4972 4483
rect 5748 4477 5788 4483
rect 5796 4477 5852 4483
rect 5940 4477 5980 4483
rect 6132 4477 6156 4483
rect 20 4457 284 4463
rect 564 4457 1004 4463
rect 1012 4457 1068 4463
rect 2212 4457 2380 4463
rect 2388 4457 2492 4463
rect 2516 4457 2716 4463
rect 2756 4457 2892 4463
rect 2900 4457 3004 4463
rect 3316 4457 3372 4463
rect 3444 4457 3500 4463
rect 3604 4457 3740 4463
rect 4132 4457 4284 4463
rect 4292 4457 4348 4463
rect 4500 4457 4508 4463
rect 4516 4457 4556 4463
rect 116 4437 684 4443
rect 916 4437 1324 4443
rect 1668 4437 1820 4443
rect 1828 4437 1964 4443
rect 1972 4437 1980 4443
rect 2260 4437 2492 4443
rect 2756 4437 3084 4443
rect 3092 4437 3180 4443
rect 3236 4437 3468 4443
rect 3924 4437 3996 4443
rect 4004 4437 4076 4443
rect 4196 4437 4204 4443
rect 4468 4437 4524 4443
rect 5716 4437 6028 4443
rect 6132 4437 6252 4443
rect 6285 4437 6291 4443
rect 2276 4417 2684 4423
rect 2724 4417 2956 4423
rect 3076 4417 3356 4423
rect 3444 4417 3548 4423
rect 4420 4417 4540 4423
rect 5716 4417 6172 4423
rect 1560 4414 1608 4416
rect 1560 4406 1564 4414
rect 1574 4406 1580 4414
rect 1588 4406 1594 4414
rect 1604 4406 1608 4414
rect 1560 4404 1608 4406
rect 4632 4414 4680 4416
rect 4632 4406 4636 4414
rect 4646 4406 4652 4414
rect 4660 4406 4666 4414
rect 4676 4406 4680 4414
rect 4632 4404 4680 4406
rect 244 4397 828 4403
rect 852 4397 1180 4403
rect 2356 4397 2460 4403
rect 2884 4397 3196 4403
rect 3876 4397 3932 4403
rect 5540 4397 6252 4403
rect -19 4377 44 4383
rect 52 4377 268 4383
rect 1012 4377 1212 4383
rect 1220 4377 1260 4383
rect 1412 4377 1468 4383
rect 1492 4377 1532 4383
rect 1540 4377 1660 4383
rect 1988 4377 2012 4383
rect 2020 4377 2092 4383
rect 2100 4377 2396 4383
rect 3188 4377 3260 4383
rect 3380 4377 3580 4383
rect 5748 4377 6156 4383
rect 580 4357 684 4363
rect 996 4357 1036 4363
rect 1428 4357 1644 4363
rect 1972 4357 1996 4363
rect 2004 4357 2076 4363
rect 2084 4357 2572 4363
rect 3172 4357 3356 4363
rect 3364 4357 3404 4363
rect 5588 4357 5916 4363
rect 5988 4357 6012 4363
rect 6036 4357 6188 4363
rect 6212 4357 6291 4363
rect -19 4337 12 4343
rect 20 4337 44 4343
rect 388 4337 412 4343
rect 420 4337 476 4343
rect 580 4337 604 4343
rect 1012 4337 1116 4343
rect 1348 4337 1388 4343
rect 1684 4337 1724 4343
rect 2052 4337 2140 4343
rect 2436 4337 2508 4343
rect 2596 4337 2636 4343
rect 2644 4337 2668 4343
rect 3348 4337 3388 4343
rect 3444 4337 3452 4343
rect 3700 4337 3820 4343
rect 4004 4337 4044 4343
rect 4052 4337 4108 4343
rect 5060 4337 5084 4343
rect 5172 4337 5244 4343
rect 5444 4337 5580 4343
rect 5620 4337 5804 4343
rect 5828 4337 5996 4343
rect 6068 4337 6092 4343
rect 6116 4337 6227 4343
rect 180 4317 220 4323
rect 436 4317 700 4323
rect 708 4317 748 4323
rect 756 4317 812 4323
rect 1140 4317 1164 4323
rect 1428 4317 1516 4323
rect 1572 4317 1660 4323
rect 1700 4317 1804 4323
rect 2196 4317 2284 4323
rect 2292 4317 2300 4323
rect 2404 4317 2444 4323
rect 2452 4317 2732 4323
rect 3012 4317 3052 4323
rect 3060 4317 3164 4323
rect 3172 4317 3228 4323
rect 3428 4317 3500 4323
rect 4212 4317 4284 4323
rect 4388 4317 4444 4323
rect 4852 4317 4876 4323
rect 5140 4317 5244 4323
rect 5284 4317 5356 4323
rect 5604 4317 5740 4323
rect 5821 4317 6012 4323
rect -19 4297 -13 4303
rect 68 4297 220 4303
rect 228 4297 316 4303
rect 468 4297 604 4303
rect 612 4297 716 4303
rect 740 4297 796 4303
rect 1140 4297 1244 4303
rect 1252 4297 1276 4303
rect 1412 4297 1452 4303
rect 1508 4297 1740 4303
rect 2228 4297 2268 4303
rect 2404 4297 2556 4303
rect 2564 4297 2604 4303
rect 2756 4297 2812 4303
rect 2964 4297 3180 4303
rect 3268 4297 3276 4303
rect 3396 4297 3436 4303
rect 3492 4297 3660 4303
rect 3668 4297 3676 4303
rect 3684 4297 3724 4303
rect 3748 4297 3772 4303
rect 3940 4297 4060 4303
rect 4068 4297 4124 4303
rect 4228 4297 4364 4303
rect 4692 4297 5116 4303
rect 5124 4297 5164 4303
rect 5300 4297 5628 4303
rect 5636 4297 5644 4303
rect 5684 4297 5724 4303
rect 5748 4297 5804 4303
rect 52 4277 92 4283
rect 116 4277 140 4283
rect 148 4277 172 4283
rect 340 4277 348 4283
rect 452 4277 508 4283
rect 788 4277 940 4283
rect 964 4277 1020 4283
rect 1236 4277 1308 4283
rect 1364 4277 1500 4283
rect 1508 4277 1708 4283
rect 1716 4277 1756 4283
rect 1972 4277 2364 4283
rect 2372 4277 2412 4283
rect 2420 4277 2460 4283
rect 2740 4277 2764 4283
rect 2900 4277 3036 4283
rect 3044 4277 3148 4283
rect 3156 4277 3212 4283
rect 3412 4277 3452 4283
rect 3732 4277 3788 4283
rect 3812 4277 3884 4283
rect 3892 4277 3932 4283
rect 4436 4277 4460 4283
rect 4468 4277 4492 4283
rect 4932 4277 4988 4283
rect 5236 4277 5276 4283
rect 5284 4277 5331 4283
rect 372 4257 636 4263
rect 692 4257 748 4263
rect 788 4257 828 4263
rect 1540 4257 1644 4263
rect 1876 4257 1996 4263
rect 2212 4257 2220 4263
rect 2308 4257 2540 4263
rect 2548 4257 2620 4263
rect 2676 4257 2684 4263
rect 3524 4257 3564 4263
rect 3572 4257 3580 4263
rect 3636 4257 3724 4263
rect 3732 4257 3820 4263
rect 4084 4257 4140 4263
rect 4148 4257 4172 4263
rect 4468 4257 4588 4263
rect 4612 4257 4844 4263
rect 4900 4257 4940 4263
rect 5300 4257 5308 4263
rect 5325 4263 5331 4277
rect 5556 4277 5580 4283
rect 5620 4277 5660 4283
rect 5821 4283 5827 4317
rect 6068 4317 6140 4323
rect 6148 4317 6204 4323
rect 6221 4323 6227 4337
rect 6221 4317 6291 4323
rect 5844 4297 5868 4303
rect 5924 4297 5996 4303
rect 6004 4297 6092 4303
rect 5821 4277 5836 4283
rect 5892 4277 5932 4283
rect 6020 4277 6044 4283
rect 6132 4277 6140 4283
rect 5325 4257 5740 4263
rect 5853 4263 5859 4276
rect 5844 4257 5859 4263
rect 5940 4257 5964 4263
rect 6036 4257 6092 4263
rect 276 4237 364 4243
rect 468 4237 556 4243
rect 772 4237 812 4243
rect 852 4237 1052 4243
rect 1124 4237 1196 4243
rect 1204 4237 1420 4243
rect 2036 4237 2268 4243
rect 2276 4237 2332 4243
rect 3252 4237 3420 4243
rect 3428 4237 3532 4243
rect 3716 4237 3852 4243
rect 3860 4237 3900 4243
rect 4052 4237 4140 4243
rect 4564 4237 4588 4243
rect 4884 4237 4956 4243
rect 5284 4237 5532 4243
rect 5588 4237 5628 4243
rect 5668 4237 5708 4243
rect 5748 4237 5852 4243
rect 5956 4237 6060 4243
rect 6132 4237 6156 4243
rect 6221 4243 6227 4296
rect 6285 4263 6291 4283
rect 6269 4257 6291 4263
rect 6221 4237 6236 4243
rect -19 4217 -13 4223
rect 596 4217 876 4223
rect 884 4217 972 4223
rect 1044 4217 1324 4223
rect 1332 4217 1484 4223
rect 1492 4217 1548 4223
rect 1860 4217 1916 4223
rect 1924 4217 2028 4223
rect 2100 4217 2364 4223
rect 3540 4217 3644 4223
rect 4180 4217 5244 4223
rect 5412 4217 5596 4223
rect 5716 4217 5740 4223
rect 5796 4217 5900 4223
rect 6269 4223 6275 4257
rect 6285 4237 6291 4243
rect 6052 4217 6275 4223
rect 3112 4214 3160 4216
rect 3112 4206 3116 4214
rect 3126 4206 3132 4214
rect 3140 4206 3146 4214
rect 3156 4206 3160 4214
rect 3112 4204 3160 4206
rect 500 4197 860 4203
rect 868 4197 956 4203
rect 1060 4197 1132 4203
rect 1444 4197 1580 4203
rect 1588 4197 1740 4203
rect 2116 4197 2220 4203
rect 2228 4197 2460 4203
rect 2580 4197 2732 4203
rect 2836 4197 2860 4203
rect 2868 4197 2924 4203
rect 2932 4197 2972 4203
rect 3316 4197 3564 4203
rect 4244 4197 4732 4203
rect 4756 4197 5164 4203
rect 5236 4197 5388 4203
rect 5460 4197 5564 4203
rect 5581 4197 5843 4203
rect 692 4177 732 4183
rect 1076 4177 1276 4183
rect 1565 4177 1708 4183
rect 1565 4164 1571 4177
rect 1956 4177 2044 4183
rect 2052 4177 2268 4183
rect 2388 4177 2540 4183
rect 2564 4177 2748 4183
rect 2756 4177 2796 4183
rect 3140 4177 3276 4183
rect 3508 4177 3548 4183
rect 3556 4177 3564 4183
rect 3572 4177 3612 4183
rect 4580 4177 4604 4183
rect 4852 4177 5100 4183
rect 5108 4177 5164 4183
rect 5581 4183 5587 4197
rect 5428 4177 5587 4183
rect 5652 4177 5820 4183
rect 5837 4183 5843 4197
rect 5972 4197 6188 4203
rect 5837 4177 6067 4183
rect 548 4157 604 4163
rect 612 4157 652 4163
rect 660 4157 684 4163
rect 804 4157 892 4163
rect 932 4157 1164 4163
rect 1300 4157 1356 4163
rect 1412 4157 1564 4163
rect 1700 4157 1884 4163
rect 1892 4157 1948 4163
rect 2116 4157 2252 4163
rect 2285 4157 2380 4163
rect 2285 4144 2291 4157
rect 2388 4157 2412 4163
rect 2484 4157 2556 4163
rect 2708 4157 2812 4163
rect 2820 4157 2956 4163
rect 3364 4157 3516 4163
rect 3556 4157 3772 4163
rect 4068 4157 4124 4163
rect 4468 4157 4524 4163
rect 4564 4157 4828 4163
rect 5012 4157 5107 4163
rect 5101 4144 5107 4157
rect 5156 4157 5244 4163
rect 5252 4157 5308 4163
rect 5364 4157 5404 4163
rect 5636 4157 5676 4163
rect 5700 4157 5724 4163
rect 5732 4157 5756 4163
rect 5789 4157 6044 4163
rect 116 4137 220 4143
rect 340 4137 396 4143
rect 532 4137 588 4143
rect 740 4137 844 4143
rect 852 4137 1132 4143
rect 1140 4137 1164 4143
rect 1364 4137 1628 4143
rect 1636 4137 1820 4143
rect 2020 4137 2044 4143
rect 2164 4137 2236 4143
rect 2324 4137 2396 4143
rect 2404 4137 2508 4143
rect 3092 4137 3219 4143
rect 20 4117 124 4123
rect 276 4117 812 4123
rect 909 4117 940 4123
rect 909 4104 915 4117
rect 1140 4117 1164 4123
rect 1220 4117 1292 4123
rect 1332 4117 1676 4123
rect 1684 4117 1868 4123
rect 1876 4117 1916 4123
rect 2004 4117 2060 4123
rect 2084 4117 2156 4123
rect 2308 4117 2428 4123
rect 2660 4117 2684 4123
rect 2948 4117 3196 4123
rect 3213 4123 3219 4137
rect 3236 4137 3308 4143
rect 3316 4137 3372 4143
rect 3396 4137 3436 4143
rect 3444 4137 3548 4143
rect 3636 4137 3740 4143
rect 3748 4137 3820 4143
rect 3988 4137 4108 4143
rect 4228 4137 4284 4143
rect 4388 4137 4780 4143
rect 4964 4137 5036 4143
rect 5108 4137 5180 4143
rect 5364 4137 5676 4143
rect 5684 4137 5708 4143
rect 5789 4143 5795 4157
rect 6061 4163 6067 4177
rect 6100 4177 6204 4183
rect 6061 4157 6108 4163
rect 6132 4157 6163 4163
rect 5741 4137 5795 4143
rect 3213 4117 3628 4123
rect 3636 4117 3660 4123
rect 3796 4117 3996 4123
rect 4212 4117 4332 4123
rect 4340 4117 4412 4123
rect 4452 4117 4876 4123
rect 4916 4117 4924 4123
rect 4932 4117 5036 4123
rect 5060 4117 5155 4123
rect -19 4097 236 4103
rect 372 4097 380 4103
rect 500 4097 620 4103
rect 836 4097 844 4103
rect 868 4097 908 4103
rect 948 4097 1244 4103
rect 1316 4097 1356 4103
rect 1396 4097 2316 4103
rect 2580 4097 2652 4103
rect 2660 4097 2668 4103
rect 2820 4097 2892 4103
rect 2948 4097 2956 4103
rect 3012 4097 3180 4103
rect 3188 4097 3244 4103
rect 4116 4097 4140 4103
rect 4148 4097 4172 4103
rect 4260 4097 4268 4103
rect 4340 4097 4348 4103
rect 4436 4097 4492 4103
rect 4500 4097 4604 4103
rect 4772 4097 4940 4103
rect 4948 4097 4988 4103
rect 5149 4103 5155 4117
rect 5252 4117 5324 4123
rect 5741 4123 5747 4137
rect 5844 4137 6012 4143
rect 6157 4143 6163 4157
rect 6180 4157 6252 4163
rect 6132 4137 6147 4143
rect 6157 4137 6195 4143
rect 5652 4117 5747 4123
rect 5764 4117 6028 4123
rect 6141 4123 6147 4137
rect 6141 4117 6172 4123
rect 5149 4097 5244 4103
rect 5293 4097 5420 4103
rect 244 4077 700 4083
rect 836 4077 1228 4083
rect 1268 4077 1516 4083
rect 1668 4077 1836 4083
rect 1988 4077 2204 4083
rect 2212 4077 2252 4083
rect 2644 4077 2700 4083
rect 2884 4077 3100 4083
rect 3284 4077 3372 4083
rect 3748 4077 3804 4083
rect 3812 4077 3980 4083
rect 4148 4077 4316 4083
rect 4324 4077 4396 4083
rect 4468 4077 4476 4083
rect 4628 4077 4668 4083
rect 4708 4077 4844 4083
rect 5293 4083 5299 4097
rect 5604 4097 5628 4103
rect 5652 4097 5660 4103
rect 5796 4097 5836 4103
rect 5869 4097 6083 4103
rect 4964 4077 5299 4083
rect 5364 4077 5388 4083
rect 5396 4077 5420 4083
rect 5668 4077 5676 4083
rect 5869 4083 5875 4097
rect 5700 4077 5875 4083
rect 5892 4077 5948 4083
rect 6077 4083 6083 4097
rect 6189 4103 6195 4137
rect 6180 4097 6195 4103
rect 6260 4097 6291 4103
rect 6077 4077 6220 4083
rect 196 4057 284 4063
rect 452 4057 588 4063
rect 852 4057 1084 4063
rect 1092 4057 1116 4063
rect 1204 4057 1468 4063
rect 1476 4057 1580 4063
rect 1588 4057 1804 4063
rect 2116 4057 2188 4063
rect 2196 4057 2236 4063
rect 2468 4057 2604 4063
rect 2708 4057 2780 4063
rect 3060 4057 3404 4063
rect 3412 4057 3596 4063
rect 3812 4057 4076 4063
rect 4132 4057 4748 4063
rect 4916 4057 5020 4063
rect 5028 4057 5052 4063
rect 5060 4057 5116 4063
rect 5172 4057 5260 4063
rect 5412 4057 5436 4063
rect 5492 4057 5676 4063
rect 5684 4057 5724 4063
rect 5876 4057 5964 4063
rect 6068 4057 6092 4063
rect 6164 4057 6188 4063
rect 436 4037 588 4043
rect 804 4037 1036 4043
rect 1092 4037 2076 4043
rect 2084 4037 2124 4043
rect 2132 4037 2156 4043
rect 2276 4037 2332 4043
rect 2340 4037 2636 4043
rect 2660 4037 2892 4043
rect 2980 4037 3068 4043
rect 3172 4037 3468 4043
rect 4404 4037 4780 4043
rect 4884 4037 4972 4043
rect 4980 4037 5004 4043
rect 5396 4037 5516 4043
rect 5684 4037 5868 4043
rect 5924 4037 6188 4043
rect 84 4017 332 4023
rect 340 4017 492 4023
rect 724 4017 1052 4023
rect 1060 4017 1100 4023
rect 1844 4017 2220 4023
rect 2932 4017 3324 4023
rect 3428 4017 3532 4023
rect 5012 4017 5100 4023
rect 5300 4017 5452 4023
rect 5908 4017 6108 4023
rect 6116 4017 6140 4023
rect 1560 4014 1608 4016
rect 1560 4006 1564 4014
rect 1574 4006 1580 4014
rect 1588 4006 1594 4014
rect 1604 4006 1608 4014
rect 1560 4004 1608 4006
rect 4632 4014 4680 4016
rect 4632 4006 4636 4014
rect 4646 4006 4652 4014
rect 4660 4006 4666 4014
rect 4676 4006 4680 4014
rect 4632 4004 4680 4006
rect 180 3997 332 4003
rect 708 3997 1404 4003
rect 1972 3997 1996 4003
rect 2036 3997 2220 4003
rect 3892 3997 4124 4003
rect 4756 3997 5772 4003
rect 5828 3997 5884 4003
rect 5908 3997 5932 4003
rect 5956 3997 5980 4003
rect 6132 3997 6236 4003
rect -19 3977 -13 3983
rect 676 3977 1100 3983
rect 1428 3977 1484 3983
rect 1508 3977 1644 3983
rect 2036 3977 2236 3983
rect 3348 3977 3580 3983
rect 3588 3977 3676 3983
rect 3700 3977 3980 3983
rect 3988 3977 4092 3983
rect 4324 3977 4588 3983
rect 4445 3964 4451 3977
rect 4788 3977 4892 3983
rect 5812 3977 5868 3983
rect 5876 3977 6028 3983
rect 20 3957 588 3963
rect 596 3957 908 3963
rect 1044 3957 1196 3963
rect 1284 3957 1436 3963
rect 1924 3957 2204 3963
rect 3428 3957 3740 3963
rect 3748 3957 3788 3963
rect 3956 3957 4012 3963
rect 4020 3957 4044 3963
rect 4068 3957 4300 3963
rect 4308 3957 4364 3963
rect 5092 3957 5196 3963
rect 5364 3957 5916 3963
rect 5988 3957 6028 3963
rect 6036 3957 6076 3963
rect 6148 3957 6172 3963
rect 132 3937 204 3943
rect 372 3937 556 3943
rect 708 3937 732 3943
rect 804 3937 876 3943
rect 948 3937 972 3943
rect 1156 3937 1468 3943
rect 2148 3937 2332 3943
rect 2564 3937 2604 3943
rect 2612 3937 2748 3943
rect 2852 3937 3388 3943
rect 3396 3937 3404 3943
rect 3412 3937 3468 3943
rect 3492 3937 3596 3943
rect 3604 3937 3660 3943
rect 3924 3937 4188 3943
rect 4196 3937 4252 3943
rect 4340 3937 4428 3943
rect 5508 3937 5580 3943
rect 5588 3937 5740 3943
rect 5844 3937 5884 3943
rect 5940 3937 6060 3943
rect 6068 3937 6252 3943
rect 6285 3937 6291 3943
rect -19 3917 -13 3923
rect 276 3917 412 3923
rect 836 3917 892 3923
rect 916 3917 1052 3923
rect 1060 3917 1180 3923
rect 1188 3917 1420 3923
rect 1908 3917 2044 3923
rect 2548 3917 2572 3923
rect 2580 3917 2620 3923
rect 2628 3917 2716 3923
rect 2788 3917 2828 3923
rect 2964 3917 3052 3923
rect 3076 3917 3148 3923
rect 3204 3917 3276 3923
rect 3556 3917 3724 3923
rect 3732 3917 3772 3923
rect 3908 3917 4044 3923
rect 4084 3917 4156 3923
rect 4180 3917 4220 3923
rect 4317 3917 4348 3923
rect 4317 3904 4323 3917
rect 4468 3917 4588 3923
rect 4596 3917 4700 3923
rect 4724 3917 4828 3923
rect 5220 3917 5244 3923
rect 5380 3917 5516 3923
rect 5524 3917 5660 3923
rect 5716 3917 6124 3923
rect 6132 3917 6172 3923
rect 116 3897 236 3903
rect 244 3897 364 3903
rect 404 3897 476 3903
rect 660 3897 796 3903
rect 820 3897 947 3903
rect 941 3884 947 3897
rect 964 3897 1068 3903
rect 1108 3897 1452 3903
rect 1460 3897 1660 3903
rect 1876 3897 1964 3903
rect 1972 3897 1996 3903
rect 2724 3897 2764 3903
rect 2980 3897 3036 3903
rect 3188 3897 3244 3903
rect 3252 3897 3340 3903
rect 3412 3897 3436 3903
rect 3492 3897 3516 3903
rect 3636 3897 3852 3903
rect 3988 3897 4060 3903
rect 4068 3897 4092 3903
rect 4116 3897 4236 3903
rect 4276 3897 4316 3903
rect 4340 3897 4396 3903
rect 4516 3897 4588 3903
rect 5012 3897 5084 3903
rect 5108 3897 5148 3903
rect 5172 3897 5196 3903
rect 5204 3897 5260 3903
rect 5572 3897 5660 3903
rect 5828 3897 5884 3903
rect 5901 3897 6220 3903
rect -19 3877 12 3883
rect 180 3877 252 3883
rect 644 3877 652 3883
rect 660 3877 908 3883
rect 948 3877 1020 3883
rect 1044 3877 1132 3883
rect 1204 3877 1292 3883
rect 1348 3877 1516 3883
rect 1620 3877 2060 3883
rect 2260 3877 2396 3883
rect 2404 3877 2636 3883
rect 2660 3877 2748 3883
rect 2756 3877 2812 3883
rect 3012 3877 3308 3883
rect 3332 3877 3564 3883
rect 3844 3877 3900 3883
rect 4052 3877 4236 3883
rect 4276 3877 4316 3883
rect 4836 3877 4860 3883
rect 4900 3877 5004 3883
rect 5140 3877 5292 3883
rect 5300 3877 5388 3883
rect 5540 3877 5644 3883
rect 5652 3877 5708 3883
rect 5901 3883 5907 3897
rect 5732 3877 5907 3883
rect 5972 3877 6044 3883
rect 6132 3877 6156 3883
rect 260 3857 348 3863
rect 644 3857 668 3863
rect 692 3857 1100 3863
rect 1108 3857 1372 3863
rect 1396 3857 1452 3863
rect 1460 3857 1820 3863
rect 1844 3857 1868 3863
rect 1892 3857 1932 3863
rect 1988 3857 2268 3863
rect 2276 3857 2380 3863
rect 2516 3857 2780 3863
rect 3220 3857 3555 3863
rect 20 3837 44 3843
rect 244 3837 412 3843
rect 676 3837 700 3843
rect 756 3837 844 3843
rect 1124 3837 1132 3843
rect 1140 3837 1196 3843
rect 1220 3837 1740 3843
rect 1844 3837 1852 3843
rect 2180 3837 2300 3843
rect 2308 3837 2588 3843
rect 2612 3837 2716 3843
rect 2756 3837 2828 3843
rect 2836 3837 2892 3843
rect 2932 3837 3180 3843
rect 3188 3837 3276 3843
rect 3284 3837 3436 3843
rect 3549 3843 3555 3857
rect 3572 3857 3580 3863
rect 3860 3857 3916 3863
rect 4292 3857 4588 3863
rect 4964 3857 5020 3863
rect 5076 3857 5100 3863
rect 5108 3857 5548 3863
rect 5700 3857 5852 3863
rect 5908 3857 5932 3863
rect 5956 3857 5980 3863
rect 6036 3857 6124 3863
rect 6148 3857 6172 3863
rect 3549 3837 3596 3843
rect 3604 3837 3708 3843
rect 3716 3837 4012 3843
rect 4612 3837 4732 3843
rect 5060 3837 5132 3843
rect 5252 3837 5276 3843
rect 5300 3837 5356 3843
rect 5364 3837 5948 3843
rect 6020 3837 6156 3843
rect 132 3817 172 3823
rect 340 3817 412 3823
rect 452 3817 540 3823
rect 628 3817 636 3823
rect 708 3817 860 3823
rect 964 3817 1324 3823
rect 1412 3817 1580 3823
rect 1636 3817 1708 3823
rect 1796 3817 1820 3823
rect 2260 3817 2396 3823
rect 2516 3817 2764 3823
rect 2772 3817 3084 3823
rect 3204 3817 3244 3823
rect 3284 3817 3356 3823
rect 3380 3817 3420 3823
rect 3428 3817 3452 3823
rect 3508 3817 3612 3823
rect 3700 3817 3756 3823
rect 3764 3817 3820 3823
rect 3908 3817 3964 3823
rect 4164 3817 4188 3823
rect 4404 3817 4428 3823
rect 4532 3817 4652 3823
rect 4660 3817 4844 3823
rect 4852 3817 5500 3823
rect 5517 3817 5724 3823
rect 3112 3814 3160 3816
rect 3112 3806 3116 3814
rect 3126 3806 3132 3814
rect 3140 3806 3146 3814
rect 3156 3806 3160 3814
rect 3112 3804 3160 3806
rect 228 3797 380 3803
rect 612 3797 764 3803
rect 772 3797 796 3803
rect 820 3797 972 3803
rect 1028 3797 1212 3803
rect 1412 3797 1484 3803
rect 1780 3797 2124 3803
rect 2132 3797 2188 3803
rect 2388 3797 2572 3803
rect 2612 3797 2668 3803
rect 2676 3797 2844 3803
rect 2852 3797 2892 3803
rect 3060 3797 3084 3803
rect 3828 3797 3852 3803
rect 4404 3797 4540 3803
rect 4564 3797 4604 3803
rect 4612 3797 4780 3803
rect 5517 3803 5523 3817
rect 5828 3817 6076 3823
rect 5140 3797 5523 3803
rect 5668 3797 5692 3803
rect 5780 3797 5820 3803
rect 5940 3797 5964 3803
rect 5988 3797 6124 3803
rect 6196 3797 6243 3803
rect -19 3777 -13 3783
rect 548 3777 684 3783
rect 852 3777 860 3783
rect 900 3777 1004 3783
rect 1012 3777 1116 3783
rect 1156 3777 1420 3783
rect 1716 3777 1852 3783
rect 1860 3777 1884 3783
rect 2500 3777 2828 3783
rect 2916 3777 2956 3783
rect 2964 3777 3308 3783
rect 3316 3777 3324 3783
rect 3348 3777 3548 3783
rect 3572 3777 3596 3783
rect 4244 3777 4284 3783
rect 4500 3777 4700 3783
rect 4724 3777 4796 3783
rect 5284 3777 5292 3783
rect 5316 3777 5372 3783
rect 5524 3777 5596 3783
rect 5652 3777 5660 3783
rect 5924 3777 5964 3783
rect 5972 3777 6156 3783
rect 6196 3777 6220 3783
rect 404 3757 460 3763
rect 660 3757 732 3763
rect 740 3757 780 3763
rect 964 3757 1052 3763
rect 1380 3757 1436 3763
rect 1940 3757 1996 3763
rect 2052 3757 2284 3763
rect 2292 3757 2348 3763
rect 2484 3757 2508 3763
rect 2644 3757 2764 3763
rect 3060 3757 3340 3763
rect 3444 3757 3628 3763
rect 4084 3757 4156 3763
rect 4484 3757 4508 3763
rect 4644 3757 4892 3763
rect 5556 3757 5612 3763
rect 5716 3757 5772 3763
rect 5812 3757 5868 3763
rect 5956 3757 5980 3763
rect 6052 3757 6140 3763
rect 6237 3763 6243 3797
rect 6228 3757 6243 3763
rect 6253 3763 6259 3776
rect 6253 3757 6275 3763
rect 148 3737 172 3743
rect 180 3737 188 3743
rect 308 3737 476 3743
rect 516 3737 572 3743
rect 580 3737 908 3743
rect 1108 3737 1164 3743
rect 1300 3737 1548 3743
rect 1988 3737 2060 3743
rect 2068 3737 2092 3743
rect 2516 3737 2572 3743
rect 2612 3737 2652 3743
rect 2932 3737 2972 3743
rect 3012 3737 3084 3743
rect 3092 3737 3180 3743
rect 3364 3737 3500 3743
rect 3540 3737 3612 3743
rect 3668 3737 3708 3743
rect 3764 3737 3788 3743
rect 3956 3737 4012 3743
rect 4228 3737 4252 3743
rect 4820 3737 4860 3743
rect 4916 3737 4940 3743
rect 4948 3737 5052 3743
rect 5092 3737 5116 3743
rect 5204 3737 5260 3743
rect 5428 3737 5452 3743
rect 5476 3737 5596 3743
rect 5636 3737 5708 3743
rect 5764 3737 5804 3743
rect 5828 3737 6028 3743
rect 6196 3737 6220 3743
rect 6244 3737 6252 3743
rect 84 3717 108 3723
rect 244 3717 316 3723
rect 484 3717 716 3723
rect 740 3717 828 3723
rect 852 3717 1356 3723
rect 1364 3717 1388 3723
rect 1396 3717 1436 3723
rect 1460 3717 1532 3723
rect 1556 3717 1756 3723
rect 1780 3717 1820 3723
rect 1828 3717 1868 3723
rect 1956 3717 2012 3723
rect 2100 3717 2140 3723
rect 2148 3717 2204 3723
rect 2276 3717 2444 3723
rect 2468 3717 2748 3723
rect 3060 3717 3068 3723
rect 3076 3717 3212 3723
rect 3220 3717 3596 3723
rect 4004 3717 4076 3723
rect 4116 3717 4332 3723
rect 4340 3717 4412 3723
rect 4724 3717 4956 3723
rect 5412 3717 5516 3723
rect 5588 3717 5756 3723
rect 5796 3717 5884 3723
rect 6093 3717 6124 3723
rect 20 3697 124 3703
rect 132 3697 172 3703
rect 180 3697 220 3703
rect 340 3697 412 3703
rect 468 3697 492 3703
rect 788 3697 812 3703
rect 820 3697 844 3703
rect 884 3697 940 3703
rect 964 3697 1020 3703
rect 1140 3697 1164 3703
rect 1332 3697 1500 3703
rect 1620 3697 1676 3703
rect 2269 3697 2332 3703
rect 2269 3684 2275 3697
rect 2372 3697 2492 3703
rect 2820 3697 2924 3703
rect 3284 3697 3340 3703
rect 3348 3697 3468 3703
rect 3492 3697 3532 3703
rect 3556 3697 3676 3703
rect 3732 3697 3772 3703
rect 4052 3697 4076 3703
rect 4164 3697 4300 3703
rect 4340 3697 4396 3703
rect 5229 3703 5235 3716
rect 5229 3697 5644 3703
rect 5812 3697 5900 3703
rect 6093 3703 6099 3717
rect 6164 3717 6236 3723
rect 5940 3697 6099 3703
rect 6116 3697 6172 3703
rect 6269 3703 6275 3757
rect 6228 3697 6275 3703
rect -19 3677 -13 3683
rect 52 3677 268 3683
rect 372 3677 604 3683
rect 788 3677 956 3683
rect 1252 3677 1356 3683
rect 1396 3677 1420 3683
rect 1444 3677 1644 3683
rect 2116 3677 2268 3683
rect 2324 3677 2396 3683
rect 2532 3677 2588 3683
rect 3012 3677 3084 3683
rect 3124 3677 3308 3683
rect 3508 3677 3580 3683
rect 4100 3677 4140 3683
rect 4148 3677 4204 3683
rect 5028 3677 5436 3683
rect 5460 3677 5788 3683
rect 5956 3677 5996 3683
rect 6004 3677 6028 3683
rect 6109 3677 6124 3683
rect 372 3657 412 3663
rect 484 3657 524 3663
rect 804 3657 860 3663
rect 1172 3657 1228 3663
rect 1236 3657 1468 3663
rect 1652 3657 1660 3663
rect 2052 3657 2412 3663
rect 2420 3657 2732 3663
rect 4196 3657 4204 3663
rect 4212 3657 4236 3663
rect 4644 3657 4748 3663
rect 4756 3657 5164 3663
rect 5453 3663 5459 3676
rect 5188 3657 5459 3663
rect 5636 3657 5676 3663
rect 5684 3657 5820 3663
rect 5860 3657 6076 3663
rect 6109 3663 6115 3677
rect 6084 3657 6115 3663
rect 6132 3657 6220 3663
rect 308 3637 444 3643
rect 580 3637 716 3643
rect 900 3637 940 3643
rect 1188 3637 1308 3643
rect 1316 3637 1436 3643
rect 1460 3637 1804 3643
rect 1812 3637 1836 3643
rect 1844 3637 1884 3643
rect 1940 3637 2380 3643
rect 2388 3637 2524 3643
rect 2804 3637 2860 3643
rect 2868 3637 2876 3643
rect 3124 3637 3404 3643
rect 3412 3637 3436 3643
rect 3508 3637 3836 3643
rect 4212 3637 4364 3643
rect 4468 3637 4908 3643
rect 4916 3637 5084 3643
rect 5396 3637 5420 3643
rect 5492 3637 5532 3643
rect 5540 3637 5868 3643
rect 5940 3637 6092 3643
rect 6100 3637 6124 3643
rect 6148 3637 6188 3643
rect -19 3617 -13 3623
rect 372 3617 428 3623
rect 1140 3617 1260 3623
rect 2372 3617 2428 3623
rect 2484 3617 2652 3623
rect 2756 3617 3004 3623
rect 3044 3617 3228 3623
rect 3348 3617 3532 3623
rect 4708 3617 5340 3623
rect 5492 3617 5516 3623
rect 5533 3617 5996 3623
rect 1560 3614 1608 3616
rect 1560 3606 1564 3614
rect 1574 3606 1580 3614
rect 1588 3606 1594 3614
rect 1604 3606 1608 3614
rect 1560 3604 1608 3606
rect 4632 3614 4680 3616
rect 4632 3606 4636 3614
rect 4646 3606 4652 3614
rect 4660 3606 4666 3614
rect 4676 3606 4680 3614
rect 4632 3604 4680 3606
rect 196 3597 268 3603
rect 292 3597 332 3603
rect 404 3597 476 3603
rect 500 3597 1196 3603
rect 1284 3597 1532 3603
rect 1716 3597 1788 3603
rect 1812 3597 2012 3603
rect 2356 3597 2588 3603
rect 3284 3597 3356 3603
rect 3780 3597 3836 3603
rect 4836 3597 5116 3603
rect 5533 3603 5539 3617
rect 6116 3617 6188 3623
rect 5364 3597 5539 3603
rect 5620 3597 5772 3603
rect 5796 3597 5836 3603
rect 5924 3597 6012 3603
rect 6228 3597 6252 3603
rect 356 3577 556 3583
rect 644 3577 892 3583
rect 900 3577 908 3583
rect 932 3577 972 3583
rect 1284 3577 1980 3583
rect 2308 3577 2508 3583
rect 2516 3577 2556 3583
rect 2612 3577 2972 3583
rect 3332 3577 3628 3583
rect 3972 3577 4332 3583
rect 4596 3577 4684 3583
rect 5204 3577 5724 3583
rect 5796 3577 5948 3583
rect 6068 3577 6140 3583
rect -19 3557 -13 3563
rect 372 3557 460 3563
rect 484 3557 556 3563
rect 580 3557 716 3563
rect 788 3557 1260 3563
rect 1268 3557 1292 3563
rect 1300 3557 1340 3563
rect 1364 3557 1500 3563
rect 1540 3557 1644 3563
rect 1748 3557 1804 3563
rect 2196 3557 2236 3563
rect 2324 3557 2716 3563
rect 2724 3557 2988 3563
rect 2996 3557 3036 3563
rect 3060 3557 3468 3563
rect 3748 3557 3932 3563
rect 4068 3557 4140 3563
rect 4180 3557 4364 3563
rect 4372 3557 4444 3563
rect 4580 3557 4828 3563
rect 5524 3557 5660 3563
rect 5748 3557 5964 3563
rect 5988 3557 6131 3563
rect 6125 3544 6131 3557
rect 148 3537 268 3543
rect 468 3537 652 3543
rect 836 3537 940 3543
rect 964 3537 1244 3543
rect 1252 3537 1308 3543
rect 1364 3537 1564 3543
rect 1620 3537 2188 3543
rect 2196 3537 2284 3543
rect 2292 3537 2348 3543
rect 2628 3537 2652 3543
rect 2772 3537 2924 3543
rect 2948 3537 2956 3543
rect 3204 3537 3244 3543
rect 3316 3537 3404 3543
rect 3492 3537 3596 3543
rect 3700 3537 3724 3543
rect 4308 3537 4412 3543
rect 4420 3537 4476 3543
rect 4548 3537 4812 3543
rect 5204 3537 5228 3543
rect 5236 3537 5276 3543
rect 5460 3537 5603 3543
rect 5597 3524 5603 3537
rect 5764 3537 5820 3543
rect 5940 3537 5996 3543
rect 6052 3537 6060 3543
rect 6228 3537 6259 3543
rect -19 3517 252 3523
rect 260 3517 620 3523
rect 1076 3517 1212 3523
rect 1236 3517 1404 3523
rect 1428 3517 1580 3523
rect 1636 3517 1644 3523
rect 1700 3517 1788 3523
rect 1972 3517 2076 3523
rect 2084 3517 2172 3523
rect 2260 3517 2476 3523
rect 2500 3517 2700 3523
rect 2740 3517 2780 3523
rect 3028 3517 3212 3523
rect 3252 3517 3292 3523
rect 3364 3517 3452 3523
rect 3460 3517 3564 3523
rect 3700 3517 3724 3523
rect 4084 3517 4156 3523
rect 4276 3517 4748 3523
rect 4772 3517 4924 3523
rect 5220 3517 5404 3523
rect 5412 3517 5468 3523
rect 5604 3517 5692 3523
rect 5748 3517 5788 3523
rect 5860 3517 5900 3523
rect 6180 3517 6220 3523
rect 148 3497 156 3503
rect 164 3497 172 3503
rect 388 3497 428 3503
rect 468 3497 588 3503
rect 660 3497 860 3503
rect 868 3497 924 3503
rect 1124 3497 1180 3503
rect 1316 3497 1356 3503
rect 1396 3497 1436 3503
rect 1604 3497 1843 3503
rect 276 3477 492 3483
rect 532 3477 812 3483
rect 884 3477 1052 3483
rect 1060 3477 1164 3483
rect 1188 3477 1484 3483
rect 1588 3477 1740 3483
rect 1780 3477 1820 3483
rect 1837 3483 1843 3497
rect 1860 3497 2204 3503
rect 2212 3497 2300 3503
rect 2340 3497 2364 3503
rect 2420 3497 2684 3503
rect 2692 3497 2748 3503
rect 2980 3497 3020 3503
rect 3268 3497 3292 3503
rect 3332 3497 3532 3503
rect 3540 3497 3548 3503
rect 3748 3497 3868 3503
rect 4212 3497 4300 3503
rect 4500 3497 4924 3503
rect 4996 3497 5036 3503
rect 5044 3497 5084 3503
rect 5252 3497 5308 3503
rect 5332 3497 5436 3503
rect 5508 3497 5532 3503
rect 5556 3497 5900 3503
rect 5917 3497 5932 3503
rect 1837 3477 1948 3483
rect 1972 3477 1980 3483
rect 2036 3477 2092 3483
rect 2148 3477 2220 3483
rect 2308 3477 2348 3483
rect 2420 3477 2476 3483
rect 2500 3477 2780 3483
rect 2948 3477 3004 3483
rect 3028 3477 3116 3483
rect 3220 3477 3388 3483
rect 3412 3477 3484 3483
rect 3508 3477 3516 3483
rect 3636 3477 3660 3483
rect 3668 3477 3756 3483
rect 4164 3477 4396 3483
rect 4404 3477 4460 3483
rect 4516 3477 4540 3483
rect 4580 3477 4764 3483
rect 4820 3477 4844 3483
rect 4996 3477 5196 3483
rect 5268 3477 5564 3483
rect 5572 3477 5772 3483
rect 5917 3483 5923 3497
rect 5780 3477 5923 3483
rect 5997 3483 6003 3496
rect 6061 3483 6067 3496
rect 5940 3477 6003 3483
rect 6029 3477 6067 3483
rect 436 3457 476 3463
rect 548 3457 732 3463
rect 740 3457 844 3463
rect 996 3457 1100 3463
rect 1108 3457 1420 3463
rect 1453 3457 1692 3463
rect -19 3437 12 3443
rect 20 3437 716 3443
rect 756 3437 796 3443
rect 820 3437 1196 3443
rect 1453 3443 1459 3457
rect 1716 3457 1772 3463
rect 1796 3457 2444 3463
rect 2452 3457 2460 3463
rect 2708 3457 2796 3463
rect 2900 3457 3084 3463
rect 3348 3457 3516 3463
rect 3524 3457 3548 3463
rect 3684 3457 3852 3463
rect 3972 3457 4108 3463
rect 4148 3457 4348 3463
rect 4356 3457 4380 3463
rect 5220 3457 5244 3463
rect 5252 3457 5292 3463
rect 5444 3457 5532 3463
rect 5700 3457 5788 3463
rect 6029 3463 6035 3477
rect 5844 3457 6035 3463
rect 6109 3463 6115 3516
rect 6132 3497 6188 3503
rect 6253 3484 6259 3537
rect 6180 3477 6220 3483
rect 6285 3483 6291 3503
rect 6269 3477 6291 3483
rect 6068 3457 6099 3463
rect 6109 3457 6188 3463
rect 1220 3437 1459 3443
rect 1604 3437 1852 3443
rect 1876 3437 2252 3443
rect 2276 3437 2588 3443
rect 2676 3437 2892 3443
rect 2932 3437 2940 3443
rect 2964 3437 2988 3443
rect 2996 3437 3132 3443
rect 3284 3437 3612 3443
rect 3620 3437 3740 3443
rect 3876 3437 4012 3443
rect 4020 3437 4124 3443
rect 4260 3437 5004 3443
rect 5268 3437 5292 3443
rect 5332 3437 5372 3443
rect 5540 3437 5852 3443
rect 5860 3437 5948 3443
rect 5988 3437 6076 3443
rect 6093 3443 6099 3457
rect 6269 3463 6275 3477
rect 6228 3457 6275 3463
rect 6285 3457 6291 3463
rect 6093 3437 6108 3443
rect 356 3417 380 3423
rect 420 3417 460 3423
rect 468 3417 524 3423
rect 724 3417 748 3423
rect 868 3417 940 3423
rect 980 3417 1052 3423
rect 1156 3417 1276 3423
rect 1316 3417 1340 3423
rect 1348 3417 1372 3423
rect 1588 3417 1612 3423
rect 1620 3417 1660 3423
rect 2164 3417 2332 3423
rect 2372 3417 2604 3423
rect 3220 3417 3244 3423
rect 3268 3417 3324 3423
rect 3348 3417 3644 3423
rect 3684 3417 3836 3423
rect 3844 3417 3996 3423
rect 4468 3417 4844 3423
rect 4852 3417 4908 3423
rect 5124 3417 5164 3423
rect 5412 3417 5740 3423
rect 5796 3417 5884 3423
rect 6036 3417 6124 3423
rect 6285 3417 6291 3423
rect 3112 3414 3160 3416
rect 3112 3406 3116 3414
rect 3126 3406 3132 3414
rect 3140 3406 3146 3414
rect 3156 3406 3160 3414
rect 3112 3404 3160 3406
rect -19 3397 236 3403
rect 612 3397 668 3403
rect 708 3397 748 3403
rect 900 3397 1132 3403
rect 1284 3397 1388 3403
rect 1476 3397 1484 3403
rect 1524 3397 1932 3403
rect 2196 3397 2236 3403
rect 2429 3397 2524 3403
rect 308 3377 332 3383
rect 372 3377 444 3383
rect 708 3377 1036 3383
rect 1133 3383 1139 3396
rect 1133 3377 1308 3383
rect 1332 3377 1596 3383
rect 1684 3377 1740 3383
rect 2429 3383 2435 3397
rect 2532 3397 2636 3403
rect 2772 3397 2828 3403
rect 2836 3397 2956 3403
rect 3181 3397 3756 3403
rect 2308 3377 2435 3383
rect 2452 3377 2492 3383
rect 2516 3377 2572 3383
rect 2580 3377 2860 3383
rect 3181 3383 3187 3397
rect 3764 3397 3772 3403
rect 3828 3397 3900 3403
rect 4052 3397 4204 3403
rect 4212 3397 4412 3403
rect 4564 3397 4620 3403
rect 5636 3397 5756 3403
rect 5844 3397 6060 3403
rect 6148 3397 6204 3403
rect 2980 3377 3187 3383
rect 3204 3377 3436 3383
rect 3444 3377 3452 3383
rect 3524 3377 3628 3383
rect 3668 3377 3692 3383
rect 3764 3377 3852 3383
rect 3860 3377 4220 3383
rect 4228 3377 4284 3383
rect 4868 3377 5004 3383
rect 5012 3377 5052 3383
rect 5652 3377 5676 3383
rect 5956 3377 5996 3383
rect 6004 3377 6220 3383
rect 6285 3377 6291 3383
rect 125 3363 131 3376
rect -19 3357 172 3363
rect 292 3357 540 3363
rect 596 3357 684 3363
rect 868 3357 876 3363
rect 916 3357 1036 3363
rect 1044 3357 1052 3363
rect 1124 3357 1164 3363
rect 1380 3357 1452 3363
rect 1460 3357 1612 3363
rect 1620 3357 1676 3363
rect 1876 3357 1980 3363
rect 2372 3357 2428 3363
rect 2436 3357 2540 3363
rect 2564 3357 2748 3363
rect 2756 3357 2812 3363
rect 2836 3357 2844 3363
rect 3236 3357 3356 3363
rect 3380 3357 3420 3363
rect 3460 3357 3564 3363
rect 3572 3357 3660 3363
rect 4228 3357 4268 3363
rect 4724 3357 4828 3363
rect 4884 3357 4924 3363
rect 5076 3357 5100 3363
rect 5364 3357 5548 3363
rect 5636 3357 5660 3363
rect 5924 3357 6124 3363
rect 6180 3357 6220 3363
rect 164 3337 220 3343
rect 244 3337 284 3343
rect 292 3337 348 3343
rect 356 3337 412 3343
rect 500 3337 588 3343
rect 596 3337 604 3343
rect 628 3337 652 3343
rect 724 3337 876 3343
rect 916 3337 1244 3343
rect 1252 3337 1292 3343
rect 1444 3337 1548 3343
rect 1652 3337 1724 3343
rect 1732 3337 1788 3343
rect 2045 3337 2156 3343
rect 260 3317 828 3323
rect 845 3317 1004 3323
rect -19 3297 44 3303
rect 308 3297 316 3303
rect 532 3297 604 3303
rect 845 3303 851 3317
rect 1012 3317 1036 3323
rect 1076 3317 1100 3323
rect 1108 3317 1340 3323
rect 1412 3317 1452 3323
rect 1469 3317 1484 3323
rect 676 3297 851 3303
rect 996 3297 1084 3303
rect 1236 3297 1276 3303
rect 1332 3297 1388 3303
rect 1469 3303 1475 3317
rect 1549 3323 1555 3336
rect 2045 3324 2051 3337
rect 2292 3337 2716 3343
rect 2804 3337 2876 3343
rect 2884 3337 2908 3343
rect 3156 3337 3260 3343
rect 3364 3337 3708 3343
rect 3716 3337 4108 3343
rect 4276 3337 4396 3343
rect 4404 3337 4492 3343
rect 4612 3337 4732 3343
rect 4868 3337 4892 3343
rect 4948 3337 4972 3343
rect 5028 3337 5052 3343
rect 5460 3337 5516 3343
rect 5620 3337 5644 3343
rect 5652 3337 5708 3343
rect 5748 3337 5820 3343
rect 5860 3337 5884 3343
rect 5908 3337 5932 3343
rect 5972 3337 6012 3343
rect 6020 3337 6291 3343
rect 1549 3317 1644 3323
rect 1748 3317 1804 3323
rect 1924 3317 2044 3323
rect 2100 3317 2124 3323
rect 2228 3317 2492 3323
rect 2500 3317 2540 3323
rect 2628 3317 2652 3323
rect 2660 3317 2707 3323
rect 2701 3304 2707 3317
rect 2852 3317 2924 3323
rect 3188 3317 3228 3323
rect 3268 3317 3308 3323
rect 3316 3317 3404 3323
rect 3428 3317 3484 3323
rect 3524 3317 3532 3323
rect 3572 3317 3724 3323
rect 3940 3317 3996 3323
rect 4004 3317 4060 3323
rect 4116 3317 4236 3323
rect 4500 3317 4556 3323
rect 4852 3317 5228 3323
rect 5444 3317 5500 3323
rect 5524 3317 5580 3323
rect 5588 3317 5644 3323
rect 5716 3317 5900 3323
rect 5972 3317 6124 3323
rect 6196 3317 6236 3323
rect 1444 3297 1475 3303
rect 1892 3297 1964 3303
rect 2132 3297 2188 3303
rect 2388 3297 2444 3303
rect 2500 3297 2636 3303
rect 2644 3297 2668 3303
rect 2708 3297 3020 3303
rect 3172 3297 3324 3303
rect 3588 3297 3628 3303
rect 3636 3297 3692 3303
rect 3700 3297 3852 3303
rect 3988 3297 4028 3303
rect 4900 3297 4908 3303
rect 4916 3297 5292 3303
rect 5332 3297 5340 3303
rect 5348 3297 5452 3303
rect 5588 3297 5980 3303
rect 212 3277 268 3283
rect 276 3277 476 3283
rect 532 3277 588 3283
rect 612 3277 620 3283
rect 644 3277 716 3283
rect 724 3277 764 3283
rect 836 3277 940 3283
rect 1028 3277 1180 3283
rect 1380 3277 1644 3283
rect 1812 3277 2060 3283
rect 2068 3277 2108 3283
rect 2212 3277 2348 3283
rect 2436 3277 2476 3283
rect 2484 3277 2524 3283
rect 2612 3277 2780 3283
rect 2820 3277 2828 3283
rect 2980 3277 3004 3283
rect 3012 3277 3212 3283
rect 3396 3277 3420 3283
rect 3428 3277 3596 3283
rect 3620 3277 3676 3283
rect 3732 3277 4428 3283
rect 4596 3277 4684 3283
rect 4980 3277 5212 3283
rect 5716 3277 5740 3283
rect 5764 3277 5900 3283
rect 5924 3277 5996 3283
rect 6020 3277 6060 3283
rect 52 3257 300 3263
rect 324 3257 396 3263
rect 468 3257 572 3263
rect 589 3263 595 3276
rect 589 3257 780 3263
rect 1012 3257 1580 3263
rect 1684 3257 1964 3263
rect 2276 3257 2684 3263
rect 2692 3257 2716 3263
rect 2964 3257 3036 3263
rect 3140 3257 3292 3263
rect 3300 3257 3420 3263
rect 3540 3257 3580 3263
rect 4388 3257 4924 3263
rect 5028 3257 5676 3263
rect 5684 3257 5788 3263
rect 5828 3257 5964 3263
rect 276 3237 524 3243
rect 676 3237 1244 3243
rect 1300 3237 1772 3243
rect 1780 3237 1868 3243
rect 1972 3237 2172 3243
rect 3412 3237 3964 3243
rect 3972 3237 4012 3243
rect 5108 3237 5180 3243
rect 5188 3237 5260 3243
rect 5492 3237 5740 3243
rect 5789 3243 5795 3256
rect 5789 3237 5900 3243
rect 132 3217 172 3223
rect 212 3217 332 3223
rect 420 3217 748 3223
rect 852 3217 1020 3223
rect 1236 3217 1292 3223
rect 1812 3217 2332 3223
rect 2932 3217 3388 3223
rect 3396 3217 3500 3223
rect 3508 3217 3756 3223
rect 3924 3217 4060 3223
rect 5092 3217 5420 3223
rect 5428 3217 5820 3223
rect 5924 3217 6028 3223
rect 6132 3217 6156 3223
rect 1560 3214 1608 3216
rect 1560 3206 1564 3214
rect 1574 3206 1580 3214
rect 1588 3206 1594 3214
rect 1604 3206 1608 3214
rect 1560 3204 1608 3206
rect 4632 3214 4680 3216
rect 4632 3206 4636 3214
rect 4646 3206 4652 3214
rect 4660 3206 4666 3214
rect 4676 3206 4680 3214
rect 4632 3204 4680 3206
rect 228 3197 284 3203
rect 404 3197 652 3203
rect 660 3197 732 3203
rect 740 3197 812 3203
rect 1060 3197 1068 3203
rect 1076 3197 1132 3203
rect 1188 3197 1452 3203
rect 1940 3197 2012 3203
rect 2324 3197 2348 3203
rect 2356 3197 2412 3203
rect 3220 3197 3283 3203
rect -19 3177 172 3183
rect 564 3177 1052 3183
rect 1284 3177 1500 3183
rect 1508 3177 1532 3183
rect 2212 3177 2252 3183
rect 2564 3177 2604 3183
rect 2708 3177 2860 3183
rect 3277 3183 3283 3197
rect 3444 3197 3740 3203
rect 3780 3197 3900 3203
rect 3917 3197 4076 3203
rect 3917 3184 3923 3197
rect 4084 3197 4236 3203
rect 5076 3197 5116 3203
rect 5524 3197 5548 3203
rect 5668 3197 5836 3203
rect 5972 3197 6060 3203
rect 3277 3177 3372 3183
rect 3508 3177 3548 3183
rect 3716 3177 3820 3183
rect 3876 3177 3916 3183
rect 4564 3177 4716 3183
rect 5124 3177 5164 3183
rect 5828 3177 6012 3183
rect 276 3157 332 3163
rect 660 3157 780 3163
rect 868 3157 876 3163
rect 1044 3157 1132 3163
rect 1156 3157 1340 3163
rect 1348 3157 1452 3163
rect 1460 3157 1548 3163
rect 1556 3157 1628 3163
rect 1780 3157 1852 3163
rect 2084 3157 2124 3163
rect 2612 3157 2636 3163
rect 2644 3157 2748 3163
rect 2916 3157 3068 3163
rect 3204 3157 3260 3163
rect 3380 3157 3436 3163
rect 3476 3157 3756 3163
rect 3764 3157 3852 3163
rect 3956 3157 4156 3163
rect 4164 3157 4204 3163
rect 4548 3157 4620 3163
rect 5300 3157 5612 3163
rect 5716 3157 5916 3163
rect 5988 3157 5996 3163
rect -19 3137 364 3143
rect 372 3137 380 3143
rect 388 3137 492 3143
rect 532 3137 700 3143
rect 836 3137 1308 3143
rect 1332 3137 1372 3143
rect 1396 3137 1420 3143
rect 1524 3137 1772 3143
rect 1780 3137 1836 3143
rect 1956 3137 1996 3143
rect 2004 3137 2108 3143
rect 2692 3137 2812 3143
rect 2820 3137 2860 3143
rect 2900 3137 3180 3143
rect 3236 3137 3276 3143
rect 3476 3137 3532 3143
rect 3636 3137 4028 3143
rect 4180 3137 4204 3143
rect 4548 3137 4604 3143
rect 4996 3137 5372 3143
rect 5428 3137 5644 3143
rect 5844 3137 5868 3143
rect 6020 3137 6060 3143
rect 180 3117 204 3123
rect 452 3117 716 3123
rect 788 3117 924 3123
rect 932 3117 1036 3123
rect 1092 3117 1164 3123
rect 1172 3117 1228 3123
rect 1332 3117 1420 3123
rect 1428 3117 1676 3123
rect 1844 3117 1868 3123
rect 2148 3117 2172 3123
rect 2196 3117 2220 3123
rect 2772 3117 2844 3123
rect 2964 3117 3020 3123
rect 3044 3117 3132 3123
rect 3252 3117 3340 3123
rect 3428 3117 3644 3123
rect 3652 3117 3676 3123
rect 3684 3117 3868 3123
rect 3892 3117 4012 3123
rect 4020 3117 4092 3123
rect 4164 3117 4252 3123
rect 4436 3117 4748 3123
rect 5172 3117 5324 3123
rect 5332 3117 5500 3123
rect 5540 3117 5660 3123
rect 5684 3117 5724 3123
rect 5908 3117 5996 3123
rect 6084 3117 6156 3123
rect 6244 3117 6291 3123
rect -19 3097 -13 3103
rect 420 3097 492 3103
rect 516 3097 556 3103
rect 708 3097 828 3103
rect 836 3097 892 3103
rect 1060 3097 1116 3103
rect 1188 3097 1244 3103
rect 1316 3097 1468 3103
rect 1476 3097 1564 3103
rect 1572 3097 1660 3103
rect 1748 3097 2012 3103
rect 2020 3097 2076 3103
rect 2404 3097 2460 3103
rect 2596 3097 2652 3103
rect 2836 3097 2876 3103
rect 3012 3097 3084 3103
rect 3252 3097 3308 3103
rect 3444 3097 3571 3103
rect 3565 3084 3571 3097
rect 3604 3097 3788 3103
rect 3908 3097 3996 3103
rect 4036 3097 4092 3103
rect 4132 3097 4172 3103
rect 4180 3097 4220 3103
rect 4484 3097 4572 3103
rect 4580 3097 4844 3103
rect 4868 3097 5036 3103
rect 5044 3097 5132 3103
rect 5236 3097 5468 3103
rect 5636 3097 5660 3103
rect 5716 3097 5724 3103
rect 5748 3097 5820 3103
rect 5876 3097 5964 3103
rect 5972 3097 6092 3103
rect 164 3077 236 3083
rect 532 3077 540 3083
rect 564 3077 684 3083
rect 724 3077 812 3083
rect 884 3077 940 3083
rect 980 3077 1004 3083
rect 1012 3077 1084 3083
rect 1348 3077 1724 3083
rect 1732 3077 1852 3083
rect 1860 3077 1932 3083
rect 2020 3077 2188 3083
rect 2452 3077 2540 3083
rect 2548 3077 2668 3083
rect 2676 3077 2748 3083
rect 2868 3077 2876 3083
rect 2980 3077 3020 3083
rect 3172 3077 3500 3083
rect 3572 3077 3644 3083
rect 3796 3077 3836 3083
rect 3860 3077 3900 3083
rect 4100 3077 4460 3083
rect 4532 3077 4700 3083
rect 4740 3077 4780 3083
rect 4804 3077 5164 3083
rect 5252 3077 5340 3083
rect 5460 3077 5500 3083
rect 5620 3077 5772 3083
rect 5780 3077 5804 3083
rect 5844 3077 6028 3083
rect 6164 3077 6291 3083
rect -19 3057 -13 3063
rect 148 3057 156 3063
rect 388 3057 412 3063
rect 500 3057 556 3063
rect 813 3063 819 3076
rect 813 3057 972 3063
rect 1044 3057 1068 3063
rect 1284 3057 1356 3063
rect 1396 3057 1427 3063
rect 1421 3044 1427 3057
rect 1460 3057 1500 3063
rect 1524 3057 1804 3063
rect 1844 3057 2236 3063
rect 2292 3057 2380 3063
rect 2852 3057 2892 3063
rect 2948 3057 3212 3063
rect 3428 3057 3452 3063
rect 3524 3057 3596 3063
rect 3636 3057 3772 3063
rect 3796 3057 3964 3063
rect 4084 3057 4108 3063
rect 4196 3057 4252 3063
rect 4292 3057 4380 3063
rect 4580 3057 4588 3063
rect 4644 3057 4748 3063
rect 4836 3057 4876 3063
rect 5012 3057 5068 3063
rect 5220 3057 5292 3063
rect 5572 3057 5692 3063
rect 5700 3057 5756 3063
rect 5764 3057 5772 3063
rect 5780 3057 6156 3063
rect 6180 3057 6204 3063
rect 20 3037 92 3043
rect 196 3037 252 3043
rect 484 3037 556 3043
rect 564 3037 588 3043
rect 596 3037 652 3043
rect 724 3037 860 3043
rect 1460 3037 1756 3043
rect 1764 3037 1868 3043
rect 1876 3037 1916 3043
rect 2004 3037 2044 3043
rect 2116 3037 2316 3043
rect 2820 3037 2908 3043
rect 2932 3037 3164 3043
rect 3220 3037 3356 3043
rect 3476 3037 3532 3043
rect 3572 3037 3676 3043
rect 3732 3037 3740 3043
rect 3748 3037 3868 3043
rect 3924 3037 4012 3043
rect 4052 3037 4348 3043
rect 4596 3037 4940 3043
rect 4948 3037 5180 3043
rect 5524 3037 5836 3043
rect 5892 3037 5964 3043
rect 6036 3037 6060 3043
rect 6244 3037 6291 3043
rect 52 3017 300 3023
rect 388 3017 604 3023
rect 868 3017 1212 3023
rect 1220 3017 1324 3023
rect 1684 3017 2012 3023
rect 2324 3017 2476 3023
rect 2484 3017 2508 3023
rect 2804 3017 3004 3023
rect 3396 3017 3436 3023
rect 3460 3017 3612 3023
rect 3764 3017 3948 3023
rect 3956 3017 4140 3023
rect 4628 3017 4716 3023
rect 4724 3017 4860 3023
rect 5012 3017 5164 3023
rect 5300 3017 5388 3023
rect 5412 3017 5580 3023
rect 5604 3017 5756 3023
rect 5780 3017 5788 3023
rect 5844 3017 6060 3023
rect 3112 3014 3160 3016
rect 3112 3006 3116 3014
rect 3126 3006 3132 3014
rect 3140 3006 3146 3014
rect 3156 3006 3160 3014
rect 3112 3004 3160 3006
rect 340 2997 540 3003
rect 580 2997 748 3003
rect 1172 2997 1196 3003
rect 1396 2997 1516 3003
rect 1524 2997 1580 3003
rect 1620 2997 1884 3003
rect 1940 2997 1964 3003
rect 1972 2997 2204 3003
rect 2580 2997 2620 3003
rect 2932 2997 2972 3003
rect 3044 2997 3075 3003
rect 116 2977 204 2983
rect 301 2977 588 2983
rect 301 2964 307 2977
rect 692 2977 940 2983
rect 964 2977 1164 2983
rect 1172 2977 1372 2983
rect 1492 2977 1692 2983
rect 1700 2977 1948 2983
rect 2068 2977 2092 2983
rect 2100 2977 2156 2983
rect 2164 2977 2300 2983
rect 2596 2977 2684 2983
rect 2868 2977 2908 2983
rect 2932 2977 3036 2983
rect 3069 2983 3075 2997
rect 3188 2997 3260 3003
rect 3284 2997 3404 3003
rect 3428 2997 3852 3003
rect 3924 2997 4124 3003
rect 4260 2997 4300 3003
rect 4756 2997 4924 3003
rect 5140 2997 5308 3003
rect 5373 2997 6291 3003
rect 5373 2984 5379 2997
rect 3069 2977 3100 2983
rect 3332 2977 3404 2983
rect 3524 2977 3596 2983
rect 3604 2977 3788 2983
rect 4020 2977 4476 2983
rect 4500 2977 4684 2983
rect 4788 2977 4956 2983
rect 4964 2977 5100 2983
rect 5108 2977 5372 2983
rect 5460 2977 5628 2983
rect 5636 2977 5804 2983
rect 5828 2977 5868 2983
rect 5956 2977 5996 2983
rect 6004 2977 6124 2983
rect 308 2957 348 2963
rect 404 2957 492 2963
rect 500 2957 524 2963
rect 532 2957 748 2963
rect 964 2957 1324 2963
rect 1460 2957 1788 2963
rect 1812 2957 1836 2963
rect 1844 2957 1852 2963
rect 2052 2957 2188 2963
rect 2516 2957 2572 2963
rect 2660 2957 2796 2963
rect 2868 2957 2892 2963
rect 2964 2957 2988 2963
rect 3012 2957 3196 2963
rect 3213 2963 3219 2976
rect 3213 2957 3244 2963
rect 3316 2957 3548 2963
rect 3556 2957 4028 2963
rect 4100 2957 4140 2963
rect 4484 2957 4620 2963
rect 4708 2957 4780 2963
rect 5108 2957 5212 2963
rect 5236 2957 5260 2963
rect 5332 2957 5356 2963
rect 5524 2957 5532 2963
rect 5556 2957 5644 2963
rect 5668 2957 5708 2963
rect 5764 2957 5788 2963
rect 5812 2957 5900 2963
rect 5908 2957 5932 2963
rect 5956 2957 5980 2963
rect 6285 2957 6291 2963
rect 228 2937 460 2943
rect 532 2937 556 2943
rect 564 2937 732 2943
rect 788 2937 860 2943
rect 868 2937 908 2943
rect 948 2937 988 2943
rect 996 2937 1068 2943
rect 1076 2937 1116 2943
rect 1444 2937 1516 2943
rect 1540 2937 1644 2943
rect 1652 2937 1740 2943
rect 1796 2937 2028 2943
rect 2036 2937 2124 2943
rect 2132 2937 2284 2943
rect 2740 2937 2956 2943
rect 2964 2937 3004 2943
rect 3076 2937 3148 2943
rect 3156 2937 3196 2943
rect 3220 2937 3308 2943
rect 3492 2937 3564 2943
rect 3620 2937 3692 2943
rect 3700 2937 3756 2943
rect 3844 2937 3868 2943
rect 3956 2937 4044 2943
rect 4244 2937 4348 2943
rect 4420 2937 4508 2943
rect 4516 2937 4540 2943
rect 4772 2937 5564 2943
rect 5684 2937 5724 2943
rect 5812 2937 5964 2943
rect 5988 2937 6012 2943
rect 6116 2937 6236 2943
rect 116 2917 444 2923
rect 541 2917 604 2923
rect 541 2904 547 2917
rect 660 2917 668 2923
rect 676 2917 780 2923
rect 1172 2917 1228 2923
rect 1268 2917 1388 2923
rect 1476 2917 1708 2923
rect 1716 2917 1772 2923
rect 1780 2917 1868 2923
rect 1892 2917 1980 2923
rect 2020 2917 2108 2923
rect 2276 2917 2332 2923
rect 2340 2917 2412 2923
rect 2420 2917 2540 2923
rect 2708 2917 2732 2923
rect 2756 2917 2988 2923
rect 3060 2917 3292 2923
rect 3332 2917 3356 2923
rect 3364 2917 3372 2923
rect 3380 2917 3452 2923
rect 3492 2917 3724 2923
rect 3828 2917 4092 2923
rect 4212 2917 4307 2923
rect 4301 2904 4307 2917
rect 4468 2917 4492 2923
rect 4500 2917 4556 2923
rect 4749 2917 4796 2923
rect -19 2897 12 2903
rect 180 2897 236 2903
rect 244 2897 316 2903
rect 436 2897 476 2903
rect 484 2897 540 2903
rect 564 2897 924 2903
rect 932 2897 1148 2903
rect 1236 2897 1404 2903
rect 1412 2897 1452 2903
rect 1636 2897 1804 2903
rect 1844 2897 1996 2903
rect 2116 2897 2268 2903
rect 2276 2897 2348 2903
rect 2356 2897 2396 2903
rect 2404 2897 2492 2903
rect 2708 2897 2828 2903
rect 2884 2897 2908 2903
rect 2932 2897 2988 2903
rect 3012 2897 3036 2903
rect 3092 2897 3180 2903
rect 3188 2897 3212 2903
rect 3300 2897 3452 2903
rect 3460 2897 3468 2903
rect 3524 2897 3724 2903
rect 3844 2897 3980 2903
rect 4212 2897 4220 2903
rect 4749 2903 4755 2917
rect 5044 2917 5084 2923
rect 5172 2917 5260 2923
rect 5268 2917 5356 2923
rect 5396 2917 5580 2923
rect 5588 2917 5900 2923
rect 5917 2917 5948 2923
rect 4340 2897 4755 2903
rect 4772 2897 4812 2903
rect 4836 2897 5356 2903
rect 5396 2897 5564 2903
rect 5652 2897 5708 2903
rect 5764 2897 5788 2903
rect 5917 2903 5923 2917
rect 5972 2917 5996 2923
rect 6068 2917 6076 2923
rect 6116 2917 6156 2923
rect 6196 2917 6220 2923
rect 5812 2897 5923 2903
rect 5940 2897 6124 2903
rect 180 2877 204 2883
rect 244 2877 332 2883
rect 596 2877 620 2883
rect 628 2877 716 2883
rect 948 2877 1068 2883
rect 1325 2877 1692 2883
rect 1325 2864 1331 2877
rect 1748 2877 1788 2883
rect 1940 2877 2172 2883
rect 2388 2877 2428 2883
rect 2436 2877 2460 2883
rect 2468 2877 2524 2883
rect 2676 2877 2748 2883
rect 2772 2877 3020 2883
rect 3028 2877 3068 2883
rect 3076 2877 3276 2883
rect 3284 2877 3420 2883
rect 3508 2877 3699 2883
rect 3693 2864 3699 2877
rect 3789 2877 4012 2883
rect 276 2857 412 2863
rect 436 2857 636 2863
rect 676 2857 812 2863
rect 916 2857 956 2863
rect 1028 2857 1036 2863
rect 1108 2857 1324 2863
rect 1684 2857 1724 2863
rect 1732 2857 2044 2863
rect 2148 2857 2300 2863
rect 2756 2857 2892 2863
rect 2900 2857 3052 2863
rect 3076 2857 3276 2863
rect 3284 2857 3676 2863
rect 3789 2863 3795 2877
rect 4276 2877 4412 2883
rect 4420 2877 4540 2883
rect 4564 2877 4716 2883
rect 4980 2877 5004 2883
rect 5076 2877 5420 2883
rect 5933 2883 5939 2896
rect 5549 2877 5939 2883
rect 5549 2864 5555 2877
rect 5956 2877 6060 2883
rect 6285 2883 6291 2903
rect 6132 2877 6291 2883
rect 3764 2857 3795 2863
rect 3812 2857 3868 2863
rect 3876 2857 3916 2863
rect 3940 2857 4060 2863
rect 4196 2857 4476 2863
rect 4596 2857 5468 2863
rect 5652 2857 5740 2863
rect 5812 2857 5868 2863
rect 6068 2857 6092 2863
rect 6132 2857 6156 2863
rect 244 2837 652 2843
rect 660 2837 684 2843
rect 708 2837 828 2843
rect 948 2837 1164 2843
rect 1428 2837 1708 2843
rect 1732 2837 1900 2843
rect 1908 2837 1948 2843
rect 2628 2837 2796 2843
rect 3012 2837 3084 2843
rect 3108 2837 3372 2843
rect 3412 2837 3580 2843
rect 3604 2837 3836 2843
rect 3892 2837 4428 2843
rect 4484 2837 4979 2843
rect 84 2817 92 2823
rect 100 2817 220 2823
rect 468 2817 492 2823
rect 644 2817 924 2823
rect 2452 2817 2636 2823
rect 2724 2817 2796 2823
rect 2932 2817 2956 2823
rect 2996 2817 3084 2823
rect 3124 2817 3196 2823
rect 3220 2817 3468 2823
rect 3508 2817 3516 2823
rect 3556 2817 3884 2823
rect 4180 2817 4380 2823
rect 4973 2823 4979 2837
rect 4996 2837 5020 2843
rect 5028 2837 5292 2843
rect 5469 2843 5475 2856
rect 5364 2837 5459 2843
rect 5469 2837 5612 2843
rect 4973 2817 5196 2823
rect 5220 2817 5388 2823
rect 5412 2817 5420 2823
rect 5453 2823 5459 2837
rect 5620 2837 5724 2843
rect 5764 2837 5852 2843
rect 5876 2837 5964 2843
rect 5988 2837 6220 2843
rect 5453 2817 5548 2823
rect 5604 2817 5756 2823
rect 5780 2817 5804 2823
rect 5860 2817 5948 2823
rect 6180 2817 6220 2823
rect 1560 2814 1608 2816
rect 1560 2806 1564 2814
rect 1574 2806 1580 2814
rect 1588 2806 1594 2814
rect 1604 2806 1608 2814
rect 1560 2804 1608 2806
rect 4632 2814 4680 2816
rect 4632 2806 4636 2814
rect 4646 2806 4652 2814
rect 4660 2806 4666 2814
rect 4676 2806 4680 2814
rect 4632 2804 4680 2806
rect 724 2797 764 2803
rect 1044 2797 1100 2803
rect 1140 2797 1260 2803
rect 1396 2797 1500 2803
rect 2772 2797 2956 2803
rect 3092 2797 3388 2803
rect 3396 2797 3532 2803
rect 3540 2797 3628 2803
rect 3636 2797 4524 2803
rect 4772 2797 5052 2803
rect 5060 2797 6124 2803
rect -19 2777 -13 2783
rect 404 2777 444 2783
rect 452 2777 700 2783
rect 884 2777 1244 2783
rect 1428 2777 1532 2783
rect 1572 2777 1756 2783
rect 1764 2777 1772 2783
rect 2660 2777 2860 2783
rect 2893 2777 3180 2783
rect 2893 2764 2899 2777
rect 3220 2777 3356 2783
rect 3380 2777 3580 2783
rect 3604 2777 3724 2783
rect 3732 2777 3948 2783
rect 4004 2777 4227 2783
rect 180 2757 428 2763
rect 484 2757 588 2763
rect 596 2757 668 2763
rect 676 2757 796 2763
rect 804 2757 1036 2763
rect 1092 2757 1644 2763
rect 2180 2757 2284 2763
rect 2292 2757 2332 2763
rect 2388 2757 2732 2763
rect 2756 2757 2892 2763
rect 3005 2757 3164 2763
rect -19 2737 108 2743
rect 516 2737 652 2743
rect 660 2737 716 2743
rect 772 2737 780 2743
rect 852 2737 908 2743
rect 980 2737 1004 2743
rect 1188 2737 1388 2743
rect 1396 2737 1404 2743
rect 1476 2737 1788 2743
rect 2004 2737 2092 2743
rect 2100 2737 2188 2743
rect 2196 2737 2220 2743
rect 2420 2737 2460 2743
rect 2468 2737 2828 2743
rect 3005 2743 3011 2757
rect 3188 2757 3228 2763
rect 3476 2757 3564 2763
rect 3572 2757 3644 2763
rect 3652 2757 3740 2763
rect 3780 2757 4204 2763
rect 4221 2763 4227 2777
rect 4244 2777 4300 2783
rect 4340 2777 4428 2783
rect 4452 2777 4508 2783
rect 4868 2777 4972 2783
rect 5012 2777 5100 2783
rect 5156 2777 5180 2783
rect 5204 2777 5267 2783
rect 4221 2757 4316 2763
rect 4324 2757 4460 2763
rect 4724 2757 4892 2763
rect 4916 2757 5004 2763
rect 5140 2757 5196 2763
rect 5220 2757 5244 2763
rect 5261 2763 5267 2777
rect 5284 2777 5532 2783
rect 5540 2777 5692 2783
rect 5700 2777 5740 2783
rect 5796 2777 5820 2783
rect 5828 2777 6236 2783
rect 5261 2757 5468 2763
rect 5492 2757 5500 2763
rect 5524 2757 5996 2763
rect 6020 2757 6044 2763
rect 2868 2737 3011 2743
rect 3204 2737 3235 2743
rect 148 2717 284 2723
rect 292 2717 316 2723
rect 548 2717 604 2723
rect 660 2717 684 2723
rect 772 2717 796 2723
rect 820 2717 1052 2723
rect 1060 2717 1164 2723
rect 1213 2717 1228 2723
rect 1213 2704 1219 2717
rect 1236 2717 1516 2723
rect 1684 2717 1884 2723
rect 1972 2717 2028 2723
rect 2436 2717 2588 2723
rect 2596 2717 2620 2723
rect 2676 2717 2700 2723
rect 2804 2717 2860 2723
rect 2868 2717 2908 2723
rect 3028 2717 3084 2723
rect 3092 2717 3100 2723
rect 3172 2717 3212 2723
rect 3229 2723 3235 2737
rect 3364 2737 3404 2743
rect 3421 2737 3484 2743
rect 3421 2723 3427 2737
rect 3492 2737 3548 2743
rect 3588 2737 3628 2743
rect 3652 2737 3804 2743
rect 3828 2737 4076 2743
rect 4084 2737 4092 2743
rect 4100 2737 4124 2743
rect 4228 2737 4284 2743
rect 4308 2737 4412 2743
rect 4436 2737 5276 2743
rect 5300 2737 5731 2743
rect 5725 2724 5731 2737
rect 5748 2737 5756 2743
rect 5780 2737 5868 2743
rect 5956 2737 6012 2743
rect 6132 2737 6204 2743
rect 3229 2717 3427 2723
rect 3476 2717 3484 2723
rect 3540 2717 3660 2723
rect 3668 2717 3772 2723
rect 3780 2717 3932 2723
rect 3972 2717 4012 2723
rect 4036 2717 4044 2723
rect 4068 2717 4108 2723
rect 4157 2717 4236 2723
rect -19 2697 12 2703
rect 20 2697 60 2703
rect 68 2697 156 2703
rect 164 2697 204 2703
rect 324 2697 860 2703
rect 980 2697 1004 2703
rect 1012 2697 1212 2703
rect 1236 2697 1260 2703
rect 1268 2697 1372 2703
rect 1380 2697 1676 2703
rect 1716 2697 1740 2703
rect 1748 2697 1852 2703
rect 1860 2697 1900 2703
rect 1908 2697 1964 2703
rect 2084 2697 2108 2703
rect 2116 2697 2172 2703
rect 2180 2697 2204 2703
rect 2292 2697 2428 2703
rect 2436 2697 2476 2703
rect 2612 2697 2700 2703
rect 2836 2697 3212 2703
rect 3220 2697 3244 2703
rect 3364 2697 3628 2703
rect 3636 2697 3756 2703
rect 3780 2697 3820 2703
rect 3828 2697 3884 2703
rect 3988 2697 4044 2703
rect 4157 2703 4163 2717
rect 4308 2717 4364 2723
rect 4372 2717 4428 2723
rect 4468 2717 4524 2723
rect 4532 2717 4627 2723
rect 4100 2697 4163 2703
rect 4180 2697 4348 2703
rect 4356 2697 4412 2703
rect 4500 2697 4556 2703
rect 4596 2697 4604 2703
rect 4621 2703 4627 2717
rect 4788 2717 4796 2723
rect 4964 2717 4972 2723
rect 4980 2717 5084 2723
rect 5108 2717 5132 2723
rect 5172 2717 5244 2723
rect 5252 2717 5564 2723
rect 5572 2717 5708 2723
rect 5732 2717 5804 2723
rect 5812 2717 5836 2723
rect 5908 2717 6060 2723
rect 6068 2717 6076 2723
rect 6100 2717 6156 2723
rect 6180 2717 6220 2723
rect 4621 2697 4796 2703
rect 4820 2697 4828 2703
rect 4852 2697 5020 2703
rect 5076 2697 5564 2703
rect 5572 2697 5644 2703
rect 5652 2697 5660 2703
rect 5700 2697 5756 2703
rect 5828 2697 5900 2703
rect 6020 2697 6028 2703
rect 6036 2697 6092 2703
rect 6100 2697 6124 2703
rect 6212 2697 6291 2703
rect 52 2677 140 2683
rect 212 2677 252 2683
rect 372 2677 412 2683
rect 516 2677 588 2683
rect 596 2677 684 2683
rect 724 2677 1052 2683
rect 1108 2677 1484 2683
rect 1556 2677 1660 2683
rect 1700 2677 1708 2683
rect 1892 2677 1980 2683
rect 2260 2677 2300 2683
rect 2308 2677 2348 2683
rect 2484 2677 2732 2683
rect 2781 2683 2787 2696
rect 2756 2677 2787 2683
rect 2804 2677 2844 2683
rect 3028 2677 3212 2683
rect 3284 2677 3308 2683
rect 3316 2677 3388 2683
rect 3524 2677 3836 2683
rect 3844 2677 3916 2683
rect 3924 2677 3948 2683
rect 4404 2677 4572 2683
rect 4660 2677 4748 2683
rect 4756 2677 4812 2683
rect 4932 2677 4988 2683
rect 5060 2677 5532 2683
rect 5588 2677 5628 2683
rect 5636 2677 5692 2683
rect 5700 2677 5772 2683
rect 5828 2677 5884 2683
rect 5908 2677 5964 2683
rect 5997 2683 6003 2696
rect 5997 2677 6012 2683
rect 6036 2677 6044 2683
rect 6052 2677 6092 2683
rect 6148 2677 6172 2683
rect 100 2657 300 2663
rect 308 2657 460 2663
rect 468 2657 492 2663
rect 564 2657 620 2663
rect 724 2657 764 2663
rect 788 2657 908 2663
rect 932 2657 988 2663
rect 1076 2657 1132 2663
rect 1140 2657 1148 2663
rect 1156 2657 1228 2663
rect 1364 2657 1932 2663
rect 1940 2657 2060 2663
rect 2180 2657 2236 2663
rect 2324 2657 2380 2663
rect 2452 2657 2492 2663
rect 2692 2657 2780 2663
rect 2804 2657 3052 2663
rect 3060 2657 3500 2663
rect 3581 2657 3612 2663
rect 260 2637 284 2643
rect 292 2637 348 2643
rect 436 2637 892 2643
rect 932 2637 1388 2643
rect 1453 2637 1772 2643
rect 1453 2624 1459 2637
rect 1780 2637 1820 2643
rect 1956 2637 2268 2643
rect 2532 2637 2588 2643
rect 2660 2637 2684 2643
rect 2740 2637 2828 2643
rect 2868 2637 2940 2643
rect 2996 2637 3068 2643
rect 3085 2637 3180 2643
rect 116 2617 300 2623
rect 308 2617 508 2623
rect 612 2617 748 2623
rect 756 2617 812 2623
rect 836 2617 956 2623
rect 1012 2617 1020 2623
rect 1108 2617 1276 2623
rect 1284 2617 1388 2623
rect 1412 2617 1452 2623
rect 1508 2617 1532 2623
rect 1748 2617 2236 2623
rect 2244 2617 2396 2623
rect 2628 2617 2972 2623
rect 3085 2623 3091 2637
rect 3204 2637 3324 2643
rect 3348 2637 3372 2643
rect 3380 2637 3452 2643
rect 3581 2643 3587 2657
rect 3636 2657 3788 2663
rect 3796 2657 3836 2663
rect 3892 2657 3964 2663
rect 3972 2657 4028 2663
rect 4084 2657 4108 2663
rect 4404 2657 5436 2663
rect 5444 2657 5452 2663
rect 5492 2657 5596 2663
rect 5620 2657 5740 2663
rect 5764 2657 5852 2663
rect 5940 2657 6140 2663
rect 6148 2657 6236 2663
rect 6285 2657 6291 2663
rect 3476 2637 3587 2643
rect 3597 2637 4044 2643
rect 2980 2617 3091 2623
rect 3236 2617 3276 2623
rect 3300 2617 3340 2623
rect 3364 2617 3404 2623
rect 3597 2623 3603 2637
rect 4052 2637 4092 2643
rect 4148 2637 4156 2643
rect 4164 2637 4204 2643
rect 4308 2637 4428 2643
rect 4580 2637 4876 2643
rect 4964 2637 5036 2643
rect 5124 2637 5180 2643
rect 5316 2637 5596 2643
rect 5620 2637 5660 2643
rect 5684 2637 5724 2643
rect 5748 2637 5811 2643
rect 3444 2617 3603 2623
rect 3620 2617 3708 2623
rect 3764 2617 3788 2623
rect 3828 2617 4140 2623
rect 4180 2617 5132 2623
rect 5156 2617 5212 2623
rect 5220 2617 5548 2623
rect 5588 2617 5788 2623
rect 5805 2623 5811 2637
rect 5844 2637 6028 2643
rect 6036 2637 6076 2643
rect 6148 2637 6188 2643
rect 5805 2617 5836 2623
rect 5860 2617 5900 2623
rect 5924 2617 5996 2623
rect 6164 2617 6188 2623
rect 3112 2614 3160 2616
rect 3112 2606 3116 2614
rect 3126 2606 3132 2614
rect 3140 2606 3146 2614
rect 3156 2606 3160 2614
rect 3112 2604 3160 2606
rect 612 2597 652 2603
rect 772 2597 812 2603
rect 836 2597 876 2603
rect 900 2597 940 2603
rect 948 2597 1068 2603
rect 1348 2597 1356 2603
rect 1412 2597 1884 2603
rect 1892 2597 1996 2603
rect 2708 2597 2940 2603
rect 3268 2597 3532 2603
rect 3604 2597 4188 2603
rect 4228 2597 4684 2603
rect 4724 2597 5164 2603
rect 5245 2597 5292 2603
rect 276 2577 524 2583
rect 660 2577 1196 2583
rect 1252 2577 1436 2583
rect 1444 2577 1484 2583
rect 1524 2577 1580 2583
rect 1588 2577 1804 2583
rect 1876 2577 2108 2583
rect 2116 2577 2300 2583
rect 2372 2577 2700 2583
rect 2756 2577 3139 2583
rect 340 2557 476 2563
rect 516 2557 572 2563
rect 708 2557 1052 2563
rect 1060 2557 1068 2563
rect 1108 2557 1148 2563
rect 1236 2557 1916 2563
rect 1924 2557 1948 2563
rect 2020 2557 2124 2563
rect 2132 2557 2316 2563
rect 2788 2557 2988 2563
rect 3133 2563 3139 2577
rect 3156 2577 3180 2583
rect 3268 2577 3468 2583
rect 3476 2577 3532 2583
rect 3620 2577 3692 2583
rect 3748 2577 3980 2583
rect 4052 2577 4060 2583
rect 4452 2577 4508 2583
rect 4516 2577 4844 2583
rect 5245 2583 5251 2597
rect 5412 2597 5948 2603
rect 5965 2597 6076 2603
rect 5133 2577 5251 2583
rect 3133 2557 3164 2563
rect 3188 2557 3356 2563
rect 3364 2557 3644 2563
rect 3732 2557 3884 2563
rect 3892 2557 3932 2563
rect 4276 2557 4380 2563
rect 4404 2557 4652 2563
rect 5133 2563 5139 2577
rect 5268 2577 5756 2583
rect 5965 2583 5971 2597
rect 5773 2577 5971 2583
rect 4708 2557 5139 2563
rect 5156 2557 5212 2563
rect 5236 2557 5308 2563
rect 5364 2557 5372 2563
rect 5773 2563 5779 2577
rect 6020 2577 6188 2583
rect 5444 2557 5779 2563
rect 5796 2557 5836 2563
rect 5981 2563 5987 2576
rect 5908 2557 5987 2563
rect 6036 2557 6092 2563
rect 6116 2557 6236 2563
rect 196 2537 316 2543
rect 468 2537 492 2543
rect 500 2537 508 2543
rect 532 2537 572 2543
rect 788 2537 812 2543
rect 852 2537 1132 2543
rect 1149 2543 1155 2556
rect 1149 2537 1292 2543
rect 1332 2537 1660 2543
rect 1485 2524 1491 2537
rect 1716 2537 1788 2543
rect 1949 2543 1955 2556
rect 1949 2537 2012 2543
rect 2164 2537 2380 2543
rect 2388 2537 2412 2543
rect 2516 2537 2524 2543
rect 2676 2537 2796 2543
rect 2852 2537 3260 2543
rect 3293 2537 3372 2543
rect 132 2517 140 2523
rect 244 2517 668 2523
rect 756 2517 1251 2523
rect -19 2497 12 2503
rect 20 2497 60 2503
rect 68 2497 172 2503
rect 180 2497 220 2503
rect 420 2497 444 2503
rect 516 2497 556 2503
rect 692 2497 1084 2503
rect 1108 2497 1164 2503
rect 1245 2503 1251 2517
rect 1284 2517 1468 2523
rect 1524 2517 1612 2523
rect 1700 2517 1740 2523
rect 2276 2517 2428 2523
rect 2452 2517 2508 2523
rect 2516 2517 2572 2523
rect 2580 2517 2652 2523
rect 2836 2517 2844 2523
rect 2884 2517 2924 2523
rect 2996 2517 3164 2523
rect 3293 2523 3299 2537
rect 3396 2537 3404 2543
rect 3412 2537 3420 2543
rect 3460 2537 3484 2543
rect 3540 2537 3596 2543
rect 3716 2537 3740 2543
rect 3844 2537 3964 2543
rect 4004 2537 4060 2543
rect 4212 2537 4252 2543
rect 4285 2537 4332 2543
rect 3204 2517 3299 2523
rect 3316 2517 3756 2523
rect 3796 2517 3900 2523
rect 3908 2517 3916 2523
rect 4285 2523 4291 2537
rect 4420 2537 4476 2543
rect 4484 2537 4524 2543
rect 4564 2537 4588 2543
rect 4612 2537 4812 2543
rect 4836 2537 4940 2543
rect 4948 2537 5004 2543
rect 5140 2537 5228 2543
rect 5252 2537 5260 2543
rect 5284 2537 5324 2543
rect 5332 2537 5420 2543
rect 5476 2537 5564 2543
rect 5588 2537 5676 2543
rect 5684 2537 5708 2543
rect 5716 2537 5852 2543
rect 5924 2537 6108 2543
rect 4020 2517 4291 2523
rect 4308 2517 4460 2523
rect 4596 2517 5388 2523
rect 5444 2517 5516 2523
rect 5540 2517 5596 2523
rect 5668 2517 5836 2523
rect 5844 2517 5932 2523
rect 6004 2517 6028 2523
rect 6052 2517 6124 2523
rect 6164 2517 6188 2523
rect 1245 2497 1580 2503
rect 1588 2497 1900 2503
rect 1908 2497 1980 2503
rect 1988 2497 2076 2503
rect 2228 2497 2476 2503
rect 2500 2497 2668 2503
rect 2708 2497 2908 2503
rect 2964 2497 3020 2503
rect 3252 2497 3324 2503
rect 3412 2497 3548 2503
rect 3556 2497 3676 2503
rect 3684 2497 3708 2503
rect 3732 2497 3788 2503
rect 3860 2497 4076 2503
rect 4084 2497 4124 2503
rect 4260 2497 4284 2503
rect 4292 2497 4332 2503
rect 4436 2497 4572 2503
rect 4692 2497 5116 2503
rect 5140 2497 5740 2503
rect 5812 2497 5932 2503
rect 5988 2497 6156 2503
rect 228 2477 364 2483
rect 468 2477 492 2483
rect 820 2477 860 2483
rect 980 2477 1132 2483
rect 1364 2477 1420 2483
rect 1428 2477 1516 2483
rect 1524 2477 1548 2483
rect 1700 2477 1708 2483
rect 2004 2477 2460 2483
rect 2468 2477 2556 2483
rect 2596 2477 2828 2483
rect 2925 2483 2931 2496
rect 2925 2477 2940 2483
rect 3028 2477 3212 2483
rect 3236 2477 3340 2483
rect 3348 2477 3468 2483
rect 3476 2477 3500 2483
rect 3588 2477 3820 2483
rect 3892 2477 4236 2483
rect 4244 2477 4316 2483
rect 4404 2477 4636 2483
rect 4644 2477 4828 2483
rect 4868 2477 4924 2483
rect 5108 2477 5244 2483
rect 5284 2477 5340 2483
rect 5348 2477 5468 2483
rect 5476 2477 5500 2483
rect 5524 2477 5884 2483
rect 5924 2477 5948 2483
rect 5972 2477 6204 2483
rect 404 2457 748 2463
rect 756 2457 908 2463
rect 916 2457 924 2463
rect 1012 2457 1404 2463
rect 1428 2457 1740 2463
rect 1972 2457 2124 2463
rect 2132 2457 2188 2463
rect 2340 2457 2524 2463
rect 2532 2457 2572 2463
rect 2612 2457 2716 2463
rect 2788 2457 3308 2463
rect 3380 2457 3452 2463
rect 3476 2457 3612 2463
rect 3668 2457 3724 2463
rect 3748 2457 3804 2463
rect 3828 2457 3868 2463
rect 3924 2457 4044 2463
rect 4084 2457 4268 2463
rect 4292 2457 4380 2463
rect 4925 2463 4931 2476
rect 4420 2457 5052 2463
rect 5124 2457 5548 2463
rect 5556 2457 5772 2463
rect 5796 2457 5884 2463
rect 5940 2457 6092 2463
rect 52 2437 108 2443
rect 532 2437 844 2443
rect 852 2437 1036 2443
rect 1076 2437 2252 2443
rect 2260 2437 2348 2443
rect 2372 2437 2620 2443
rect 2644 2437 2924 2443
rect 2932 2437 3068 2443
rect 3092 2437 3772 2443
rect 3805 2443 3811 2456
rect 3805 2437 3980 2443
rect 4132 2437 4172 2443
rect 4301 2437 4556 2443
rect 116 2417 140 2423
rect 308 2417 332 2423
rect 340 2417 364 2423
rect 436 2417 620 2423
rect 628 2417 1068 2423
rect 1188 2417 1228 2423
rect 1332 2417 1452 2423
rect 2004 2417 2252 2423
rect 2276 2417 2572 2423
rect 2612 2417 2956 2423
rect 2980 2417 2988 2423
rect 3012 2417 3100 2423
rect 3268 2417 3292 2423
rect 3300 2417 3436 2423
rect 3524 2417 3580 2423
rect 3732 2417 3756 2423
rect 4301 2423 4307 2437
rect 4580 2437 4748 2443
rect 4788 2437 4876 2443
rect 4884 2437 6060 2443
rect 6100 2437 6124 2443
rect 3828 2417 4307 2423
rect 4324 2417 4604 2423
rect 4772 2417 4812 2423
rect 4836 2417 5532 2423
rect 5588 2417 5923 2423
rect 1560 2414 1608 2416
rect 1560 2406 1564 2414
rect 1574 2406 1580 2414
rect 1588 2406 1594 2414
rect 1604 2406 1608 2414
rect 1560 2404 1608 2406
rect 4632 2414 4680 2416
rect 4632 2406 4636 2414
rect 4646 2406 4652 2414
rect 4660 2406 4666 2414
rect 4676 2406 4680 2414
rect 4632 2404 4680 2406
rect -19 2397 12 2403
rect 20 2397 60 2403
rect 148 2397 188 2403
rect 196 2397 396 2403
rect 964 2397 1420 2403
rect 1652 2397 1948 2403
rect 2068 2397 2172 2403
rect 2356 2397 2844 2403
rect 2900 2397 2924 2403
rect 3060 2397 3244 2403
rect 3348 2397 3468 2403
rect 3492 2397 3884 2403
rect 3956 2397 3996 2403
rect 4052 2397 4220 2403
rect 4260 2397 4556 2403
rect 4708 2397 5020 2403
rect 5124 2397 5900 2403
rect 5917 2403 5923 2417
rect 6084 2417 6140 2423
rect 5917 2397 5996 2403
rect 84 2377 108 2383
rect 164 2377 316 2383
rect 324 2377 380 2383
rect 653 2377 1388 2383
rect -19 2357 92 2363
rect 100 2357 124 2363
rect 132 2357 156 2363
rect 212 2357 236 2363
rect 260 2357 364 2363
rect 653 2363 659 2377
rect 1476 2377 1724 2383
rect 1844 2377 1996 2383
rect 2100 2377 2268 2383
rect 2484 2377 2700 2383
rect 2724 2377 3116 2383
rect 3156 2377 3404 2383
rect 3412 2377 3484 2383
rect 3620 2377 3820 2383
rect 3844 2377 4172 2383
rect 4180 2377 4204 2383
rect 4212 2377 4364 2383
rect 4388 2377 4444 2383
rect 4500 2377 4588 2383
rect 4660 2377 4716 2383
rect 4788 2377 4828 2383
rect 4884 2377 4940 2383
rect 4964 2377 4972 2383
rect 4980 2377 4988 2383
rect 5108 2377 5260 2383
rect 5284 2377 5388 2383
rect 5460 2377 5580 2383
rect 5668 2377 5804 2383
rect 6004 2377 6156 2383
rect 372 2357 659 2363
rect 676 2357 1676 2363
rect 1732 2357 1772 2363
rect 1780 2357 1852 2363
rect 1860 2357 1900 2363
rect 1988 2357 2204 2363
rect 2516 2357 3132 2363
rect 3348 2357 3452 2363
rect 3469 2357 4172 2363
rect 3469 2344 3475 2357
rect 4180 2357 5420 2363
rect 5556 2357 5804 2363
rect 5812 2357 5852 2363
rect 5876 2357 6012 2363
rect 6164 2357 6188 2363
rect 6244 2357 6259 2363
rect 276 2337 348 2343
rect 356 2337 412 2343
rect 452 2337 476 2343
rect 628 2337 636 2343
rect 660 2337 1676 2343
rect 1684 2337 1804 2343
rect 1812 2337 1836 2343
rect 1908 2337 2140 2343
rect 2324 2337 2396 2343
rect 2404 2337 2460 2343
rect 2580 2337 2636 2343
rect 2676 2337 3468 2343
rect 3492 2337 3612 2343
rect 3652 2337 3756 2343
rect 3780 2337 3820 2343
rect 3924 2337 4604 2343
rect 4612 2337 4908 2343
rect 5044 2337 5100 2343
rect 5188 2337 5276 2343
rect 5332 2337 5404 2343
rect 5748 2337 5996 2343
rect 6116 2337 6236 2343
rect 6253 2343 6259 2357
rect 6253 2337 6307 2343
rect -19 2317 12 2323
rect 20 2317 284 2323
rect 292 2317 444 2323
rect 452 2317 556 2323
rect 596 2317 668 2323
rect 756 2317 828 2323
rect 868 2317 988 2323
rect 996 2317 1068 2323
rect 1108 2317 1132 2323
rect 1220 2317 1276 2323
rect 1316 2317 1356 2323
rect 1364 2317 1372 2323
rect 1444 2317 1740 2323
rect 1748 2317 1820 2323
rect 1892 2317 1932 2323
rect 1956 2317 2012 2323
rect 2052 2317 2291 2323
rect 196 2297 220 2303
rect 244 2297 348 2303
rect 356 2297 428 2303
rect 468 2297 572 2303
rect 676 2297 700 2303
rect 724 2297 748 2303
rect 836 2297 892 2303
rect 916 2297 940 2303
rect 948 2297 1020 2303
rect 1044 2297 1084 2303
rect 1204 2297 1292 2303
rect 1348 2297 1452 2303
rect 1508 2297 1516 2303
rect 1540 2297 1564 2303
rect 2205 2297 2268 2303
rect 2205 2284 2211 2297
rect 2285 2303 2291 2317
rect 2420 2317 2476 2323
rect 2484 2317 2796 2323
rect 2820 2317 2892 2323
rect 2909 2317 2956 2323
rect 2285 2297 2508 2303
rect 2564 2297 2620 2303
rect 2660 2297 2684 2303
rect 2708 2297 2764 2303
rect 2909 2303 2915 2317
rect 2980 2317 3004 2323
rect 3028 2317 3084 2323
rect 3188 2317 3212 2323
rect 3268 2317 3292 2323
rect 3332 2317 3388 2323
rect 3444 2317 3516 2323
rect 3604 2317 3884 2323
rect 3892 2317 3900 2323
rect 3972 2317 4060 2323
rect 4068 2317 4140 2323
rect 4148 2317 4188 2323
rect 4196 2317 4348 2323
rect 4404 2317 4428 2323
rect 4500 2317 4636 2323
rect 4644 2317 4764 2323
rect 4964 2317 5084 2323
rect 5108 2317 5164 2323
rect 5172 2317 5212 2323
rect 5300 2317 5356 2323
rect 5476 2317 5484 2323
rect 5572 2317 5628 2323
rect 5636 2317 5900 2323
rect 5908 2317 5932 2323
rect 6052 2317 6108 2323
rect 2884 2297 2915 2303
rect 2948 2297 3020 2303
rect 3044 2297 3148 2303
rect 3188 2297 3196 2303
rect 3268 2297 3308 2303
rect 3316 2297 3331 2303
rect 116 2277 140 2283
rect 164 2277 540 2283
rect 708 2277 1116 2283
rect 1140 2277 1148 2283
rect 1156 2277 1420 2283
rect 1524 2277 1708 2283
rect 1796 2277 1884 2283
rect 2068 2277 2204 2283
rect 2260 2277 2316 2283
rect 2324 2277 2364 2283
rect 2420 2277 2844 2283
rect 2852 2277 2908 2283
rect 2964 2277 2988 2283
rect 3060 2277 3308 2283
rect 3325 2283 3331 2297
rect 3364 2297 3404 2303
rect 3460 2297 3500 2303
rect 3732 2297 3916 2303
rect 4276 2297 4332 2303
rect 4340 2297 4492 2303
rect 4516 2297 4588 2303
rect 4596 2297 4668 2303
rect 4756 2297 4780 2303
rect 4813 2297 5132 2303
rect 4813 2284 4819 2297
rect 5332 2297 5356 2303
rect 5668 2297 5724 2303
rect 5812 2297 5916 2303
rect 5940 2297 5996 2303
rect 3325 2277 3356 2283
rect 3492 2277 3596 2283
rect 3636 2277 3724 2283
rect 3732 2277 3964 2283
rect 3972 2277 4012 2283
rect 4436 2277 4556 2283
rect 4580 2277 4700 2283
rect 4708 2277 4764 2283
rect 4852 2277 4940 2283
rect 5012 2277 5052 2283
rect 5140 2277 5180 2283
rect 5188 2277 5292 2283
rect 5316 2277 5420 2283
rect 5444 2277 5500 2283
rect 5508 2277 5612 2283
rect 5700 2277 5868 2283
rect 5885 2277 5971 2283
rect 52 2257 268 2263
rect 308 2257 556 2263
rect 660 2257 764 2263
rect 932 2257 1036 2263
rect 1188 2257 1244 2263
rect 1252 2257 1660 2263
rect 1940 2257 2108 2263
rect 2436 2257 2508 2263
rect 2516 2257 2604 2263
rect 2676 2257 2780 2263
rect 2836 2257 3068 2263
rect 3108 2257 3164 2263
rect 3204 2257 3244 2263
rect 3284 2257 3436 2263
rect 3492 2257 3548 2263
rect 3620 2257 3859 2263
rect 52 2237 156 2243
rect 260 2237 332 2243
rect 340 2237 492 2243
rect 804 2237 828 2243
rect 836 2237 956 2243
rect 1012 2237 1068 2243
rect 1092 2237 1196 2243
rect 1380 2237 1420 2243
rect 1956 2237 2236 2243
rect 2244 2237 2252 2243
rect 2660 2237 2716 2243
rect 2724 2237 2812 2243
rect 2884 2237 2972 2243
rect 2996 2237 3084 2243
rect 3156 2237 3740 2243
rect 3764 2237 3836 2243
rect 3853 2243 3859 2257
rect 3924 2257 4092 2263
rect 4228 2257 4316 2263
rect 4548 2257 4588 2263
rect 4596 2257 4828 2263
rect 4836 2257 4956 2263
rect 4996 2257 5020 2263
rect 5028 2257 5084 2263
rect 5092 2257 5148 2263
rect 5284 2257 5468 2263
rect 5556 2257 5596 2263
rect 5885 2263 5891 2277
rect 5604 2257 5891 2263
rect 5965 2263 5971 2277
rect 6020 2277 6060 2283
rect 6084 2277 6124 2283
rect 5965 2257 6156 2263
rect 3853 2237 3996 2243
rect 4468 2237 4732 2243
rect 4756 2237 4796 2243
rect 4804 2237 4940 2243
rect 5149 2243 5155 2256
rect 5149 2237 5324 2243
rect 5652 2237 5804 2243
rect 5860 2237 5884 2243
rect 5908 2237 5932 2243
rect 5988 2237 6060 2243
rect 6100 2237 6140 2243
rect 6173 2243 6179 2296
rect 6173 2237 6188 2243
rect 84 2217 188 2223
rect 196 2217 364 2223
rect 372 2217 380 2223
rect 484 2217 540 2223
rect 964 2217 1347 2223
rect -19 2197 -13 2203
rect 212 2197 220 2203
rect 228 2197 252 2203
rect 500 2197 508 2203
rect 756 2197 844 2203
rect 868 2197 1036 2203
rect 1076 2197 1244 2203
rect 1252 2197 1276 2203
rect 1341 2203 1347 2217
rect 1364 2217 1532 2223
rect 1540 2217 1868 2223
rect 2420 2217 2492 2223
rect 2932 2217 3036 2223
rect 3188 2217 3260 2223
rect 3316 2217 3788 2223
rect 3796 2217 4028 2223
rect 4276 2217 4716 2223
rect 4772 2217 4892 2223
rect 4964 2217 5244 2223
rect 5652 2217 5708 2223
rect 5748 2217 5820 2223
rect 5828 2217 5964 2223
rect 5988 2217 6028 2223
rect 6180 2217 6252 2223
rect 3112 2214 3160 2216
rect 3112 2206 3116 2214
rect 3126 2206 3132 2214
rect 3140 2206 3146 2214
rect 3156 2206 3160 2214
rect 3112 2204 3160 2206
rect 1341 2197 1500 2203
rect 1732 2197 1996 2203
rect 2324 2197 2508 2203
rect 2573 2197 2892 2203
rect 2573 2184 2579 2197
rect 2932 2197 3036 2203
rect 3220 2197 3276 2203
rect 3380 2197 3660 2203
rect 3741 2197 4220 2203
rect 20 2177 92 2183
rect 116 2177 204 2183
rect 516 2177 876 2183
rect 1124 2177 1212 2183
rect 1412 2177 1436 2183
rect 1524 2177 2140 2183
rect 2148 2177 2172 2183
rect 2260 2177 2572 2183
rect 2884 2177 3228 2183
rect 3268 2177 3372 2183
rect 3412 2177 3516 2183
rect 3540 2177 3564 2183
rect 3741 2183 3747 2197
rect 4244 2197 4428 2203
rect 4452 2197 4499 2203
rect 3620 2177 3747 2183
rect 3860 2177 3916 2183
rect 4004 2177 4108 2183
rect 4196 2177 4220 2183
rect 4244 2177 4412 2183
rect 4420 2177 4476 2183
rect 4493 2183 4499 2197
rect 4516 2197 5148 2203
rect 5220 2197 5740 2203
rect 5764 2197 6028 2203
rect 6084 2197 6092 2203
rect 6148 2197 6156 2203
rect 4493 2177 4988 2183
rect 4996 2177 5020 2183
rect 5076 2177 5100 2183
rect 5140 2177 5324 2183
rect 5332 2177 5388 2183
rect 5716 2177 5948 2183
rect 6116 2177 6236 2183
rect 164 2157 300 2163
rect 340 2157 492 2163
rect 500 2157 588 2163
rect 596 2157 636 2163
rect 692 2157 908 2163
rect 916 2157 1004 2163
rect 1341 2157 1516 2163
rect 1341 2144 1347 2157
rect 1684 2157 2012 2163
rect 2036 2157 2092 2163
rect 2100 2157 2188 2163
rect 2308 2157 2476 2163
rect 2900 2157 2956 2163
rect 3060 2157 3068 2163
rect 3076 2157 3340 2163
rect 3412 2157 3452 2163
rect 3476 2157 3564 2163
rect 3604 2157 3740 2163
rect 3748 2157 3820 2163
rect 3908 2157 3980 2163
rect 4020 2157 4716 2163
rect 4740 2157 4844 2163
rect 4852 2157 4940 2163
rect 4980 2157 5036 2163
rect 5140 2157 5340 2163
rect 5348 2157 5404 2163
rect 5620 2157 5628 2163
rect 5956 2157 6204 2163
rect 36 2137 172 2143
rect 484 2137 652 2143
rect 884 2137 972 2143
rect 980 2137 1020 2143
rect 1044 2137 1068 2143
rect 1188 2137 1340 2143
rect 1412 2137 1820 2143
rect 1828 2137 1884 2143
rect 1908 2137 1964 2143
rect 1972 2137 2060 2143
rect 2301 2143 2307 2156
rect 2301 2137 2348 2143
rect 2580 2137 2812 2143
rect 2820 2137 2940 2143
rect 3028 2137 3052 2143
rect 3236 2137 3308 2143
rect 3348 2137 3372 2143
rect 3444 2137 3500 2143
rect 3684 2137 3708 2143
rect 3716 2137 3939 2143
rect 116 2117 140 2123
rect 244 2117 316 2123
rect 324 2117 380 2123
rect 436 2117 620 2123
rect 708 2117 780 2123
rect 1060 2117 1251 2123
rect 68 2097 108 2103
rect 468 2097 508 2103
rect 612 2097 700 2103
rect 756 2097 1180 2103
rect 1245 2103 1251 2117
rect 1268 2117 1420 2123
rect 1508 2117 1628 2123
rect 1668 2117 1708 2123
rect 2020 2117 2044 2123
rect 2132 2117 2156 2123
rect 2212 2117 2268 2123
rect 2276 2117 2364 2123
rect 2420 2117 2444 2123
rect 2596 2117 2780 2123
rect 2836 2117 3244 2123
rect 3252 2117 3420 2123
rect 3428 2117 3763 2123
rect 1245 2097 1276 2103
rect 1316 2097 1628 2103
rect 1636 2097 1756 2103
rect 1764 2097 1852 2103
rect 1908 2097 1948 2103
rect 2004 2097 2028 2103
rect 2084 2097 2252 2103
rect 2324 2097 3356 2103
rect 3364 2097 3644 2103
rect 3661 2097 3740 2103
rect 404 2077 684 2083
rect 884 2077 1260 2083
rect 1332 2077 1571 2083
rect 116 2057 140 2063
rect 308 2057 460 2063
rect 484 2057 716 2063
rect 724 2057 780 2063
rect 996 2057 1036 2063
rect 1044 2057 1100 2063
rect 1428 2057 1500 2063
rect 1565 2063 1571 2077
rect 1652 2077 1804 2083
rect 1812 2077 1868 2083
rect 1876 2077 1916 2083
rect 2260 2077 2348 2083
rect 2388 2077 2556 2083
rect 2644 2077 2732 2083
rect 2852 2077 2908 2083
rect 2964 2077 3132 2083
rect 3156 2077 3196 2083
rect 3252 2077 3292 2083
rect 3300 2077 3340 2083
rect 3412 2077 3468 2083
rect 3508 2077 3596 2083
rect 3661 2083 3667 2097
rect 3757 2103 3763 2117
rect 3780 2117 3884 2123
rect 3933 2123 3939 2137
rect 3956 2137 4028 2143
rect 4180 2137 4268 2143
rect 4308 2137 4348 2143
rect 4404 2137 4460 2143
rect 4516 2137 4604 2143
rect 4740 2137 5100 2143
rect 5156 2137 5228 2143
rect 5236 2137 5292 2143
rect 5364 2137 5628 2143
rect 5636 2137 5980 2143
rect 6004 2137 6012 2143
rect 6132 2137 6188 2143
rect 3933 2117 4012 2123
rect 4084 2117 4108 2123
rect 4212 2117 4252 2123
rect 4404 2117 4444 2123
rect 4452 2117 4524 2123
rect 4564 2117 4572 2123
rect 4580 2117 4812 2123
rect 5012 2117 5052 2123
rect 5076 2117 5132 2123
rect 5252 2117 5276 2123
rect 5357 2117 5436 2123
rect 3757 2097 3772 2103
rect 3780 2097 4844 2103
rect 5357 2103 5363 2117
rect 5444 2117 5516 2123
rect 5572 2117 5660 2123
rect 5668 2117 5724 2123
rect 5732 2117 5836 2123
rect 5940 2117 5971 2123
rect 5965 2104 5971 2117
rect 6045 2123 6051 2136
rect 6221 2124 6227 2156
rect 6020 2117 6051 2123
rect 6100 2117 6124 2123
rect 6180 2117 6204 2123
rect 4868 2097 5363 2103
rect 5396 2097 5676 2103
rect 5684 2097 5708 2103
rect 5716 2097 5772 2103
rect 5876 2097 5955 2103
rect 3613 2077 3667 2083
rect 1565 2057 1644 2063
rect 1652 2057 1724 2063
rect 1908 2057 2236 2063
rect 2436 2057 2476 2063
rect 2612 2057 2796 2063
rect 2804 2057 2844 2063
rect 2868 2057 3180 2063
rect 3204 2057 3228 2063
rect 3284 2057 3372 2063
rect 3613 2063 3619 2077
rect 3684 2077 3868 2083
rect 3908 2077 3948 2083
rect 4029 2077 4108 2083
rect 3444 2057 3619 2063
rect 3636 2057 3676 2063
rect 4029 2063 4035 2077
rect 4356 2077 4508 2083
rect 4548 2077 4588 2083
rect 4612 2077 5148 2083
rect 5156 2077 5308 2083
rect 5316 2077 5580 2083
rect 5732 2077 5868 2083
rect 5876 2077 5884 2083
rect 5949 2083 5955 2097
rect 6036 2097 6092 2103
rect 5949 2077 6044 2083
rect 6052 2077 6076 2083
rect 3748 2057 4035 2063
rect 4052 2057 4140 2063
rect 4196 2057 4540 2063
rect 4564 2057 4620 2063
rect 4628 2057 4716 2063
rect 4756 2057 4972 2063
rect 5300 2057 5484 2063
rect 5492 2057 5612 2063
rect 5652 2057 6131 2063
rect 244 2037 732 2043
rect 756 2037 940 2043
rect 1092 2037 1132 2043
rect 1300 2037 2012 2043
rect 2301 2043 2307 2056
rect 2020 2037 2396 2043
rect 2708 2037 2892 2043
rect 2900 2037 3020 2043
rect 3044 2037 3100 2043
rect 3140 2037 3580 2043
rect 3588 2037 3708 2043
rect 3716 2037 3788 2043
rect 3924 2037 4083 2043
rect 84 2017 1100 2023
rect 1124 2017 1452 2023
rect 1668 2017 1692 2023
rect 2244 2017 2332 2023
rect 2340 2017 2412 2023
rect 2452 2017 2684 2023
rect 2724 2017 3004 2023
rect 3028 2017 3100 2023
rect 3188 2017 3724 2023
rect 3732 2017 4012 2023
rect 4077 2023 4083 2037
rect 4100 2037 4284 2043
rect 4292 2037 4316 2043
rect 4324 2037 4380 2043
rect 4436 2037 4707 2043
rect 4077 2017 4348 2023
rect 4701 2023 4707 2037
rect 4724 2037 5132 2043
rect 5165 2043 5171 2056
rect 5165 2037 5356 2043
rect 5380 2037 5468 2043
rect 5508 2037 5532 2043
rect 5812 2037 6076 2043
rect 6100 2037 6108 2043
rect 6125 2043 6131 2057
rect 6125 2037 6220 2043
rect 4701 2017 4748 2023
rect 4772 2017 4956 2023
rect 4996 2017 5500 2023
rect 5540 2017 5612 2023
rect 5620 2017 5740 2023
rect 5780 2017 6028 2023
rect 6036 2017 6140 2023
rect 6301 2023 6307 2337
rect 6180 2017 6307 2023
rect 1560 2014 1608 2016
rect 1560 2006 1564 2014
rect 1574 2006 1580 2014
rect 1588 2006 1594 2014
rect 1604 2006 1608 2014
rect 1560 2004 1608 2006
rect 4632 2014 4680 2016
rect 4632 2006 4636 2014
rect 4646 2006 4652 2014
rect 4660 2006 4666 2014
rect 4676 2006 4680 2014
rect 4632 2004 4680 2006
rect 308 1997 364 2003
rect 436 1997 460 2003
rect 564 1997 588 2003
rect 884 1997 1020 2003
rect 1060 1997 1148 2003
rect 1156 1997 1228 2003
rect 1284 1997 1484 2003
rect 1652 1997 1868 2003
rect 1956 1997 2092 2003
rect 2420 1997 3532 2003
rect 3540 1997 3820 2003
rect 3828 1997 4124 2003
rect 4148 1997 4300 2003
rect 4820 1997 4828 2003
rect 4852 1997 4940 2003
rect 5908 1997 5932 2003
rect 6036 1997 6060 2003
rect 6084 1997 6236 2003
rect 404 1977 540 1983
rect 564 1977 956 1983
rect 980 1977 1356 1983
rect 1364 1977 1436 1983
rect 1652 1977 1756 1983
rect 2084 1977 2140 1983
rect 2148 1977 2492 1983
rect 2948 1977 3036 1983
rect 3076 1977 3164 1983
rect 3172 1977 3260 1983
rect 3284 1977 4108 1983
rect 4125 1983 4131 1996
rect 4125 1977 5068 1983
rect 5268 1977 5964 1983
rect 6116 1977 6124 1983
rect 212 1957 300 1963
rect 308 1957 460 1963
rect 756 1957 1164 1963
rect 1188 1957 1212 1963
rect 1220 1957 1340 1963
rect 1572 1957 1676 1963
rect 1684 1957 1724 1963
rect 2052 1957 2092 1963
rect 2100 1957 2220 1963
rect 2772 1957 2812 1963
rect 2980 1957 3180 1963
rect 3188 1957 3196 1963
rect 3220 1957 3484 1963
rect 3508 1957 3612 1963
rect 3684 1957 4044 1963
rect 4052 1957 4060 1963
rect 4420 1957 4604 1963
rect 4612 1957 4844 1963
rect 4852 1957 4876 1963
rect 4948 1957 5372 1963
rect 5428 1957 5468 1963
rect 5492 1957 5708 1963
rect 5716 1957 5852 1963
rect 5860 1957 5932 1963
rect 5956 1957 6060 1963
rect 6068 1957 6124 1963
rect 36 1937 124 1943
rect 228 1937 284 1943
rect 372 1937 380 1943
rect 484 1937 492 1943
rect 820 1937 1132 1943
rect 1140 1937 1164 1943
rect 1172 1937 1212 1943
rect 1268 1937 1324 1943
rect 1380 1937 1420 1943
rect 2093 1937 2172 1943
rect 84 1917 140 1923
rect 148 1917 572 1923
rect 596 1917 668 1923
rect 676 1917 796 1923
rect 804 1917 892 1923
rect 900 1917 908 1923
rect 964 1917 1004 1923
rect 1012 1917 1036 1923
rect 1076 1917 1100 1923
rect 1172 1917 1356 1923
rect 1380 1917 1452 1923
rect 1508 1917 1724 1923
rect 1732 1917 1804 1923
rect 1876 1917 1900 1923
rect 2093 1923 2099 1937
rect 2180 1937 2220 1943
rect 2340 1937 2348 1943
rect 2404 1937 2444 1943
rect 2516 1937 2540 1943
rect 2548 1937 2636 1943
rect 2740 1937 2764 1943
rect 2804 1937 2844 1943
rect 2877 1937 3692 1943
rect 1940 1917 2099 1923
rect 2877 1923 2883 1937
rect 3700 1937 3820 1943
rect 3828 1937 3948 1943
rect 3956 1937 5516 1943
rect 5556 1937 5692 1943
rect 5716 1937 5932 1943
rect 5940 1937 5996 1943
rect 2132 1917 2883 1923
rect 2900 1917 2956 1923
rect 2996 1917 3052 1923
rect 3108 1917 3212 1923
rect 3300 1917 3388 1923
rect 3396 1917 3516 1923
rect 3588 1917 3667 1923
rect 3661 1904 3667 1917
rect 3716 1917 3740 1923
rect 3876 1917 4236 1923
rect 4292 1917 4332 1923
rect 4356 1917 4380 1923
rect 4436 1917 4620 1923
rect 4628 1917 4828 1923
rect 4916 1917 5148 1923
rect 5156 1917 5180 1923
rect 5460 1917 5484 1923
rect 5588 1917 5644 1923
rect 5668 1917 5884 1923
rect 5892 1917 5980 1923
rect 6132 1917 6172 1923
rect 100 1897 332 1903
rect 340 1897 396 1903
rect 596 1897 636 1903
rect 644 1897 732 1903
rect 740 1897 812 1903
rect 820 1897 844 1903
rect 852 1897 876 1903
rect 948 1897 1004 1903
rect 1124 1897 1148 1903
rect 1204 1897 1292 1903
rect 1332 1897 1516 1903
rect 1524 1897 1740 1903
rect 1748 1897 1868 1903
rect 2020 1897 2060 1903
rect 2068 1897 2108 1903
rect 2196 1897 2236 1903
rect 2356 1897 2460 1903
rect 2692 1897 2748 1903
rect 2772 1897 2876 1903
rect 2980 1897 3004 1903
rect 3012 1897 3036 1903
rect 3076 1897 3100 1903
rect 3108 1897 3180 1903
rect 3284 1897 3340 1903
rect 3364 1897 3500 1903
rect 3556 1897 3644 1903
rect 3668 1897 3708 1903
rect 3748 1897 4172 1903
rect 4212 1897 4444 1903
rect 4452 1897 4492 1903
rect 4964 1897 5020 1903
rect 5140 1897 5660 1903
rect 5732 1897 5868 1903
rect 6164 1897 6172 1903
rect 6228 1897 6236 1903
rect 6285 1897 6291 1903
rect 20 1877 172 1883
rect 180 1877 476 1883
rect 484 1877 684 1883
rect 724 1877 860 1883
rect 868 1877 940 1883
rect 964 1877 1020 1883
rect 1364 1877 1436 1883
rect 1492 1877 1692 1883
rect 1732 1877 1756 1883
rect 1764 1877 1804 1883
rect 2212 1877 2268 1883
rect 2308 1877 2700 1883
rect 2868 1877 2988 1883
rect 3332 1877 3372 1883
rect 3572 1877 3788 1883
rect 3796 1877 3836 1883
rect 3940 1877 3996 1883
rect 4036 1877 4076 1883
rect 4132 1877 4204 1883
rect 4260 1877 4428 1883
rect 4468 1877 4540 1883
rect 4564 1877 4732 1883
rect 4740 1877 5244 1883
rect 5252 1877 5388 1883
rect 5405 1877 5532 1883
rect -19 1857 -13 1863
rect 68 1857 188 1863
rect 196 1857 236 1863
rect 356 1857 396 1863
rect 500 1857 732 1863
rect 868 1857 908 1863
rect 1028 1857 1116 1863
rect 1124 1857 1148 1863
rect 1284 1857 1388 1863
rect 1396 1857 1644 1863
rect 2340 1857 2348 1863
rect 2365 1857 2444 1863
rect 276 1837 348 1843
rect 372 1837 764 1843
rect 820 1837 1404 1843
rect 1492 1837 2044 1843
rect 2365 1843 2371 1857
rect 2452 1857 2588 1863
rect 2964 1857 2972 1863
rect 3044 1857 3180 1863
rect 3268 1857 3308 1863
rect 3492 1857 3548 1863
rect 3556 1857 3580 1863
rect 3604 1857 3724 1863
rect 3773 1857 3948 1863
rect 2276 1837 2371 1843
rect 2388 1837 2732 1843
rect 2932 1837 3084 1843
rect 3124 1837 3196 1843
rect 3220 1837 3452 1843
rect 3773 1843 3779 1857
rect 3988 1857 4156 1863
rect 4164 1857 4220 1863
rect 4340 1857 4476 1863
rect 4484 1857 4508 1863
rect 4532 1857 4716 1863
rect 4788 1857 4828 1863
rect 4836 1857 4860 1863
rect 5044 1857 5148 1863
rect 5188 1857 5228 1863
rect 5236 1857 5276 1863
rect 5405 1863 5411 1877
rect 5716 1877 5772 1883
rect 5876 1877 5916 1883
rect 5924 1877 5980 1883
rect 5988 1877 6028 1883
rect 6132 1877 6188 1883
rect 5364 1857 5411 1863
rect 5428 1857 5596 1863
rect 5828 1857 5884 1863
rect 6036 1857 6156 1863
rect 6196 1857 6236 1863
rect 3524 1837 3779 1843
rect 3796 1837 4188 1843
rect 4196 1837 4284 1843
rect 4292 1837 4364 1843
rect 4596 1837 4652 1843
rect 4660 1837 4748 1843
rect 4756 1837 5196 1843
rect 5220 1837 5292 1843
rect 5300 1837 5324 1843
rect 5796 1837 5964 1843
rect 6004 1837 6188 1843
rect -19 1817 -13 1823
rect 244 1817 252 1823
rect 276 1817 524 1823
rect 692 1817 844 1823
rect 852 1817 908 1823
rect 932 1817 1036 1823
rect 1076 1817 1516 1823
rect 1524 1817 1772 1823
rect 1780 1817 1820 1823
rect 2372 1817 2492 1823
rect 2500 1817 2556 1823
rect 2564 1817 2620 1823
rect 2820 1817 3068 1823
rect 3348 1817 3916 1823
rect 3924 1817 3964 1823
rect 4068 1817 4220 1823
rect 5284 1817 5372 1823
rect 5924 1817 6028 1823
rect 3112 1814 3160 1816
rect 3112 1806 3116 1814
rect 3126 1806 3132 1814
rect 3140 1806 3146 1814
rect 3156 1806 3160 1814
rect 3112 1804 3160 1806
rect 148 1797 387 1803
rect 148 1777 188 1783
rect 381 1783 387 1797
rect 429 1797 636 1803
rect 429 1783 435 1797
rect 660 1797 716 1803
rect 756 1797 940 1803
rect 1044 1797 1196 1803
rect 1204 1797 1228 1803
rect 1428 1797 1452 1803
rect 1476 1797 1628 1803
rect 2388 1797 2444 1803
rect 2452 1797 2476 1803
rect 2516 1797 2572 1803
rect 2580 1797 2636 1803
rect 2644 1797 2876 1803
rect 2900 1797 2956 1803
rect 3028 1797 3084 1803
rect 3188 1797 3356 1803
rect 3620 1797 3644 1803
rect 3892 1797 4140 1803
rect 4164 1797 4172 1803
rect 4196 1797 4364 1803
rect 4404 1797 4572 1803
rect 4724 1797 4828 1803
rect 4948 1797 5196 1803
rect 5812 1797 5820 1803
rect 381 1777 435 1783
rect 452 1777 460 1783
rect 676 1777 716 1783
rect 724 1777 796 1783
rect 804 1777 1068 1783
rect 1076 1777 1164 1783
rect 1380 1777 1388 1783
rect 1428 1777 1548 1783
rect 1684 1777 1724 1783
rect 1940 1777 1996 1783
rect 2004 1777 2060 1783
rect 2164 1777 2476 1783
rect 2804 1777 2812 1783
rect 2852 1777 2892 1783
rect 2900 1777 2940 1783
rect 2948 1777 3004 1783
rect 3124 1777 3228 1783
rect 3316 1777 3452 1783
rect 3508 1777 3596 1783
rect 3668 1777 3692 1783
rect 3828 1777 3852 1783
rect 3876 1777 4060 1783
rect 4148 1777 4316 1783
rect 4324 1777 4451 1783
rect 84 1757 380 1763
rect 388 1757 460 1763
rect 580 1757 604 1763
rect 708 1757 748 1763
rect 772 1757 828 1763
rect 836 1757 940 1763
rect 957 1757 1196 1763
rect 180 1737 236 1743
rect 356 1737 556 1743
rect 708 1737 796 1743
rect 852 1737 892 1743
rect 916 1737 924 1743
rect 957 1743 963 1757
rect 1220 1757 1260 1763
rect 1268 1757 1708 1763
rect 1780 1757 2012 1763
rect 2132 1757 2236 1763
rect 2356 1757 2604 1763
rect 2612 1757 2716 1763
rect 2740 1757 2796 1763
rect 2916 1757 3084 1763
rect 3108 1757 3196 1763
rect 3204 1757 3212 1763
rect 3229 1763 3235 1776
rect 3229 1757 3276 1763
rect 3300 1757 3388 1763
rect 3572 1757 3612 1763
rect 3636 1757 3644 1763
rect 3652 1757 3676 1763
rect 3700 1757 3708 1763
rect 3764 1757 4428 1763
rect 4445 1763 4451 1777
rect 4468 1777 4764 1783
rect 4884 1777 4988 1783
rect 4996 1777 5036 1783
rect 5348 1777 5628 1783
rect 5636 1777 5708 1783
rect 5892 1777 5996 1783
rect 6285 1777 6291 1783
rect 4445 1757 4476 1763
rect 4788 1757 4924 1763
rect 4932 1757 4972 1763
rect 4980 1757 5068 1763
rect 5268 1757 5292 1763
rect 5492 1757 5564 1763
rect 5956 1757 5971 1763
rect 932 1737 963 1743
rect 1076 1737 1244 1743
rect 1252 1737 1308 1743
rect 1316 1737 1484 1743
rect 1508 1737 1532 1743
rect 1604 1737 1692 1743
rect 1700 1737 1932 1743
rect 2068 1737 2124 1743
rect 2164 1737 2364 1743
rect 2445 1737 2588 1743
rect 196 1717 332 1723
rect 372 1717 412 1723
rect 452 1717 508 1723
rect 564 1717 636 1723
rect 660 1717 684 1723
rect 724 1717 956 1723
rect 964 1717 1004 1723
rect 1044 1717 1084 1723
rect 1140 1717 1180 1723
rect 1252 1717 1292 1723
rect 1348 1717 1468 1723
rect 1485 1723 1491 1736
rect 2445 1724 2451 1737
rect 2708 1737 2748 1743
rect 2820 1737 3020 1743
rect 3188 1737 3212 1743
rect 3220 1737 3260 1743
rect 3284 1737 3340 1743
rect 3396 1737 3660 1743
rect 3700 1737 3900 1743
rect 3908 1737 3948 1743
rect 3956 1737 4012 1743
rect 4132 1737 4396 1743
rect 4532 1737 4588 1743
rect 4804 1737 5068 1743
rect 5076 1737 5132 1743
rect 5140 1737 5308 1743
rect 5316 1737 5388 1743
rect 5396 1737 5516 1743
rect 5844 1737 5948 1743
rect 1485 1717 1868 1723
rect 1876 1717 1884 1723
rect 2116 1717 2172 1723
rect 2228 1717 2444 1723
rect 2484 1717 2604 1723
rect 2676 1717 3404 1723
rect 3412 1717 4300 1723
rect 4308 1717 4524 1723
rect 4532 1717 4684 1723
rect 4708 1717 4876 1723
rect 4900 1717 4988 1723
rect 5012 1717 5036 1723
rect 5044 1717 5308 1723
rect 5316 1717 5404 1723
rect 5428 1717 5468 1723
rect 5476 1717 5500 1723
rect 5508 1717 5596 1723
rect 5652 1717 5740 1723
rect 5965 1723 5971 1757
rect 6052 1737 6236 1743
rect 5956 1717 5971 1723
rect -19 1697 12 1703
rect 20 1697 60 1703
rect 68 1697 108 1703
rect 116 1697 156 1703
rect 420 1697 460 1703
rect 596 1697 1356 1703
rect 1380 1697 1676 1703
rect 1716 1697 1756 1703
rect 1876 1697 1932 1703
rect 2116 1697 2156 1703
rect 2196 1697 2316 1703
rect 2388 1697 2460 1703
rect 2468 1697 2524 1703
rect 2612 1697 2716 1703
rect 2724 1697 2748 1703
rect 2804 1697 3020 1703
rect 3028 1697 3228 1703
rect 3300 1697 3372 1703
rect 3556 1697 3676 1703
rect 3684 1697 3724 1703
rect 3732 1697 3916 1703
rect 4116 1697 4140 1703
rect 4244 1697 4300 1703
rect 4308 1697 4332 1703
rect 4340 1697 4572 1703
rect 4580 1697 4716 1703
rect 4740 1697 4876 1703
rect 4916 1697 5356 1703
rect 5364 1697 5372 1703
rect 5604 1697 5676 1703
rect 5684 1697 5724 1703
rect 5812 1697 5836 1703
rect 5892 1697 5980 1703
rect 6164 1697 6291 1703
rect 484 1677 860 1683
rect 1028 1677 1100 1683
rect 1108 1677 1468 1683
rect 1556 1677 1788 1683
rect 2132 1677 2156 1683
rect 2292 1677 2348 1683
rect 2356 1677 2412 1683
rect 2436 1677 2540 1683
rect 2548 1677 2572 1683
rect 2820 1677 2860 1683
rect 2932 1677 3036 1683
rect 3108 1677 3404 1683
rect 3876 1677 4092 1683
rect 4100 1677 4124 1683
rect 4276 1677 4348 1683
rect 4420 1677 5548 1683
rect 5844 1677 5868 1683
rect 6020 1677 6124 1683
rect 100 1657 876 1663
rect 900 1657 1004 1663
rect 1012 1657 1116 1663
rect 1140 1657 1164 1663
rect 1268 1657 1324 1663
rect 1364 1657 1612 1663
rect 1652 1657 1692 1663
rect 1700 1657 1836 1663
rect 1844 1657 2156 1663
rect 2164 1657 2620 1663
rect 2644 1657 2972 1663
rect 3028 1657 3436 1663
rect 3460 1657 3612 1663
rect 3629 1657 3756 1663
rect 308 1637 348 1643
rect 356 1637 492 1643
rect 516 1637 716 1643
rect 788 1637 1148 1643
rect 1156 1637 1388 1643
rect 1524 1637 1532 1643
rect 1540 1637 1852 1643
rect 2004 1637 2380 1643
rect 2404 1637 2476 1643
rect 2820 1637 3020 1643
rect 3629 1643 3635 1657
rect 3796 1657 4028 1663
rect 4212 1657 4396 1663
rect 4548 1657 4748 1663
rect 4964 1657 5084 1663
rect 5860 1657 6092 1663
rect 3204 1637 3635 1643
rect 3652 1637 3852 1643
rect 3860 1637 3932 1643
rect 4004 1637 4044 1643
rect 4052 1637 4108 1643
rect 4436 1637 4979 1643
rect 100 1617 268 1623
rect 340 1617 492 1623
rect 532 1617 588 1623
rect 660 1617 876 1623
rect 980 1617 1516 1623
rect 2052 1617 2668 1623
rect 2724 1617 2924 1623
rect 2948 1617 3228 1623
rect 3236 1617 3276 1623
rect 3469 1617 3532 1623
rect 1560 1614 1608 1616
rect 1560 1606 1564 1614
rect 1574 1606 1580 1614
rect 1588 1606 1594 1614
rect 1604 1606 1608 1614
rect 1560 1604 1608 1606
rect 52 1597 396 1603
rect 557 1597 668 1603
rect 557 1583 563 1597
rect 692 1597 732 1603
rect 829 1597 1180 1603
rect 68 1577 563 1583
rect 829 1583 835 1597
rect 1188 1597 1196 1603
rect 1284 1597 1532 1603
rect 1828 1597 2188 1603
rect 2388 1597 2844 1603
rect 3469 1603 3475 1617
rect 3556 1617 3884 1623
rect 3972 1617 4124 1623
rect 4973 1623 4979 1637
rect 4996 1637 5452 1643
rect 6052 1637 6076 1643
rect 6285 1637 6291 1643
rect 4973 1617 5148 1623
rect 5156 1617 5260 1623
rect 5476 1617 5740 1623
rect 5748 1617 5900 1623
rect 4632 1614 4680 1616
rect 4632 1606 4636 1614
rect 4646 1606 4652 1614
rect 4660 1606 4666 1614
rect 4676 1606 4680 1614
rect 4632 1604 4680 1606
rect 2884 1597 3475 1603
rect 3764 1597 3772 1603
rect 3812 1597 3932 1603
rect 3956 1597 3980 1603
rect 4084 1597 4108 1603
rect 4148 1597 4476 1603
rect 4820 1597 5036 1603
rect 5268 1597 6252 1603
rect 628 1577 835 1583
rect 932 1577 972 1583
rect 996 1577 1260 1583
rect 1348 1577 1500 1583
rect 1668 1577 2028 1583
rect 2228 1577 2268 1583
rect 2340 1577 2444 1583
rect 2468 1577 2860 1583
rect 2996 1577 3068 1583
rect 3076 1577 3212 1583
rect 3252 1577 3388 1583
rect 3460 1577 3804 1583
rect 3924 1577 4227 1583
rect 4221 1564 4227 1577
rect 4260 1577 4364 1583
rect 4372 1577 4428 1583
rect 4436 1577 4556 1583
rect 4660 1577 4956 1583
rect 5908 1577 5948 1583
rect 6212 1577 6236 1583
rect 276 1557 332 1563
rect 404 1557 428 1563
rect 436 1557 1036 1563
rect 1108 1557 1164 1563
rect 1172 1557 1292 1563
rect 1460 1557 1564 1563
rect 1700 1557 1852 1563
rect 1860 1557 1916 1563
rect 2404 1557 2732 1563
rect 2740 1557 2796 1563
rect 2932 1557 2956 1563
rect 2964 1557 2988 1563
rect 3028 1557 3068 1563
rect 3140 1557 3260 1563
rect 3316 1557 3372 1563
rect 3380 1557 3676 1563
rect 3764 1557 3852 1563
rect 3876 1557 3980 1563
rect 4068 1557 4092 1563
rect 4116 1557 4172 1563
rect 4228 1557 4268 1563
rect 4404 1557 4460 1563
rect 4820 1557 4828 1563
rect 4932 1557 5308 1563
rect 5316 1557 5356 1563
rect 5396 1557 6172 1563
rect 196 1537 412 1543
rect 420 1537 547 1543
rect -19 1517 12 1523
rect 20 1517 403 1523
rect 397 1504 403 1517
rect 436 1517 476 1523
rect 541 1523 547 1537
rect 564 1537 652 1543
rect 660 1537 812 1543
rect 916 1537 1084 1543
rect 1108 1537 1196 1543
rect 1236 1537 1292 1543
rect 1508 1537 1932 1543
rect 1940 1537 1996 1543
rect 2292 1537 2444 1543
rect 2452 1537 2700 1543
rect 2724 1537 2780 1543
rect 2836 1537 2860 1543
rect 2900 1537 2956 1543
rect 2964 1537 3244 1543
rect 3348 1537 3580 1543
rect 3732 1537 3804 1543
rect 3860 1537 4124 1543
rect 4468 1537 4908 1543
rect 4916 1537 4956 1543
rect 5108 1537 5292 1543
rect 5300 1537 5340 1543
rect 5700 1537 5836 1543
rect 5844 1537 5932 1543
rect 541 1517 588 1523
rect 676 1517 716 1523
rect 788 1517 812 1523
rect 868 1517 956 1523
rect 1044 1517 1548 1523
rect 1556 1517 1660 1523
rect 1844 1517 2060 1523
rect 2068 1517 2108 1523
rect 2180 1517 2332 1523
rect 2340 1517 2348 1523
rect 2356 1517 2380 1523
rect 2436 1517 2604 1523
rect 2637 1517 2812 1523
rect 132 1497 156 1503
rect 180 1497 204 1503
rect 212 1497 364 1503
rect 404 1497 524 1503
rect 628 1497 652 1503
rect 660 1497 1020 1503
rect 1076 1497 1100 1503
rect 1204 1497 1244 1503
rect 1316 1497 1356 1503
rect 1460 1497 1484 1503
rect 1796 1497 1836 1503
rect 1844 1497 1900 1503
rect 1924 1497 2092 1503
rect 2100 1497 2204 1503
rect 2308 1497 2364 1503
rect 2548 1497 2588 1503
rect 2637 1503 2643 1517
rect 2836 1517 3276 1523
rect 3428 1517 3468 1523
rect 3780 1517 3884 1523
rect 3908 1517 3948 1523
rect 4036 1517 4044 1523
rect 4052 1517 4236 1523
rect 4340 1517 4412 1523
rect 4500 1517 4508 1523
rect 4516 1517 4572 1523
rect 4596 1517 4764 1523
rect 4772 1517 4828 1523
rect 4980 1517 5020 1523
rect 5076 1517 5132 1523
rect 5140 1517 5164 1523
rect 5364 1517 5436 1523
rect 5732 1517 5788 1523
rect 5828 1517 5868 1523
rect 2596 1497 2643 1503
rect 2660 1497 2700 1503
rect 2772 1497 3180 1503
rect 3204 1497 3260 1503
rect 3444 1497 4108 1503
rect 4116 1497 4284 1503
rect 4292 1497 4732 1503
rect 4756 1497 4780 1503
rect 4820 1497 4860 1503
rect 4884 1497 4924 1503
rect 4948 1497 5004 1503
rect 5060 1497 5100 1503
rect 5108 1497 5196 1503
rect 5444 1497 5564 1503
rect 5700 1497 5740 1503
rect 5748 1497 5820 1503
rect 5876 1497 5948 1503
rect 20 1477 156 1483
rect 164 1477 220 1483
rect 292 1477 316 1483
rect 468 1477 508 1483
rect 580 1477 684 1483
rect 692 1477 844 1483
rect 900 1477 924 1483
rect 948 1477 988 1483
rect 1076 1477 1084 1483
rect 1140 1477 1228 1483
rect 1245 1483 1251 1496
rect 1245 1477 1724 1483
rect 1732 1477 1964 1483
rect 2164 1477 2316 1483
rect 2324 1477 2412 1483
rect 2500 1477 2556 1483
rect 2596 1477 2620 1483
rect 2660 1477 2668 1483
rect 2756 1477 3020 1483
rect 3044 1477 3132 1483
rect 3156 1477 3180 1483
rect 3284 1477 3388 1483
rect 3444 1477 3564 1483
rect 3604 1477 3660 1483
rect 3668 1477 3980 1483
rect 4036 1477 4140 1483
rect 4196 1477 4204 1483
rect 4212 1477 4252 1483
rect 4324 1477 4444 1483
rect 4468 1477 4716 1483
rect 4724 1477 4892 1483
rect 4925 1483 4931 1496
rect 4925 1477 4972 1483
rect 5428 1477 5484 1483
rect 5492 1477 5532 1483
rect 5780 1477 5788 1483
rect 5796 1477 5884 1483
rect 5924 1477 6044 1483
rect 6052 1477 6156 1483
rect 212 1457 284 1463
rect 612 1457 700 1463
rect 708 1457 732 1463
rect 772 1457 796 1463
rect 868 1457 972 1463
rect 1076 1457 1164 1463
rect 1172 1457 1212 1463
rect 1300 1457 1372 1463
rect 1588 1457 1708 1463
rect 1908 1457 1980 1463
rect 1988 1457 2012 1463
rect 2100 1457 2140 1463
rect 2196 1457 2508 1463
rect 2621 1463 2627 1476
rect 2621 1457 2716 1463
rect 2772 1457 2796 1463
rect 2884 1457 2988 1463
rect 3012 1457 3164 1463
rect 3188 1457 4284 1463
rect 4445 1463 4451 1476
rect 4445 1457 4524 1463
rect 4644 1457 4668 1463
rect 5012 1457 5052 1463
rect 5284 1457 5324 1463
rect 5332 1457 5388 1463
rect 5412 1457 5580 1463
rect 5620 1457 6028 1463
rect 596 1437 716 1443
rect 756 1437 844 1443
rect 1028 1437 1276 1443
rect 1284 1437 1660 1443
rect 2084 1437 2204 1443
rect 2244 1437 2412 1443
rect 2484 1437 2508 1443
rect 2516 1437 2684 1443
rect 2692 1437 2812 1443
rect 2820 1437 3196 1443
rect 3220 1437 3340 1443
rect 3588 1437 3644 1443
rect 3796 1437 3804 1443
rect 3876 1437 4412 1443
rect 4420 1437 4556 1443
rect 4564 1437 4796 1443
rect 4804 1437 4844 1443
rect 4996 1437 5468 1443
rect 5588 1437 5708 1443
rect 5716 1437 5772 1443
rect 6020 1437 6108 1443
rect 148 1417 348 1423
rect 532 1417 588 1423
rect 612 1417 828 1423
rect 836 1417 892 1423
rect 1060 1417 1404 1423
rect 1412 1417 1436 1423
rect 1844 1417 2492 1423
rect 2564 1417 2876 1423
rect 2932 1417 2956 1423
rect 2996 1417 3004 1423
rect 3060 1417 3084 1423
rect 3284 1417 3324 1423
rect 3412 1417 3516 1423
rect 3540 1417 3644 1423
rect 3725 1417 3916 1423
rect 3112 1414 3160 1416
rect 3112 1406 3116 1414
rect 3126 1406 3132 1414
rect 3140 1406 3146 1414
rect 3156 1406 3160 1414
rect 3112 1404 3160 1406
rect 500 1397 524 1403
rect 564 1397 748 1403
rect 884 1397 924 1403
rect 980 1397 1004 1403
rect 1012 1397 1020 1403
rect 1156 1397 1228 1403
rect 1364 1397 1420 1403
rect 2132 1397 2252 1403
rect 2260 1397 2476 1403
rect 2484 1397 2540 1403
rect 2804 1397 2812 1403
rect 2980 1397 3091 1403
rect 228 1377 252 1383
rect 260 1377 316 1383
rect 356 1377 556 1383
rect 628 1377 636 1383
rect 852 1377 908 1383
rect 932 1377 956 1383
rect 980 1377 1100 1383
rect 1204 1377 1212 1383
rect 1300 1377 1356 1383
rect 1476 1377 1628 1383
rect 1684 1377 1740 1383
rect 1972 1377 1996 1383
rect 2004 1377 2108 1383
rect 2276 1377 2316 1383
rect 2340 1377 2364 1383
rect 2708 1377 2844 1383
rect 2852 1377 2956 1383
rect 2964 1377 3036 1383
rect 3085 1383 3091 1397
rect 3188 1397 3372 1403
rect 3725 1403 3731 1417
rect 3940 1417 3948 1423
rect 4292 1417 4348 1423
rect 4356 1417 4540 1423
rect 4788 1417 5084 1423
rect 5092 1417 5180 1423
rect 5956 1417 6060 1423
rect 3428 1397 3731 1403
rect 3748 1397 4156 1403
rect 4212 1397 5132 1403
rect 5588 1397 5868 1403
rect 3085 1377 3356 1383
rect 3412 1377 3420 1383
rect 3508 1377 3532 1383
rect 3572 1377 3580 1383
rect 3636 1377 3692 1383
rect 3700 1377 3772 1383
rect 3988 1377 4316 1383
rect 4340 1377 4556 1383
rect 5764 1377 5916 1383
rect 5924 1377 5996 1383
rect 52 1357 108 1363
rect 420 1357 492 1363
rect 500 1357 620 1363
rect 628 1357 668 1363
rect 756 1357 780 1363
rect 964 1357 1580 1363
rect 1652 1357 1692 1363
rect 1716 1357 2012 1363
rect 2100 1357 2172 1363
rect 2532 1357 2659 1363
rect 212 1337 236 1343
rect 484 1337 636 1343
rect 644 1337 716 1343
rect 756 1337 780 1343
rect 820 1337 1036 1343
rect 1204 1337 1244 1343
rect 1284 1337 1340 1343
rect 1604 1337 1955 1343
rect 1949 1324 1955 1337
rect 2100 1337 2179 1343
rect 52 1317 124 1323
rect 596 1317 684 1323
rect 756 1317 924 1323
rect 996 1317 1212 1323
rect 1220 1317 1228 1323
rect 1332 1317 1532 1323
rect 1572 1317 1660 1323
rect 1668 1317 1692 1323
rect 1796 1317 1884 1323
rect 2068 1317 2140 1323
rect 2173 1323 2179 1337
rect 2196 1337 2396 1343
rect 2404 1337 2508 1343
rect 2516 1337 2556 1343
rect 2653 1343 2659 1357
rect 2676 1357 3084 1363
rect 3092 1357 3452 1363
rect 3460 1357 3628 1363
rect 3636 1357 3708 1363
rect 3924 1357 3964 1363
rect 3972 1357 4060 1363
rect 4116 1357 4140 1363
rect 4260 1357 4444 1363
rect 4452 1357 4492 1363
rect 4884 1357 4940 1363
rect 5044 1357 5196 1363
rect 5213 1357 5260 1363
rect 5213 1344 5219 1357
rect 5652 1357 5756 1363
rect 5764 1357 5852 1363
rect 2653 1337 2851 1343
rect 2173 1317 2252 1323
rect 2308 1317 2348 1323
rect 2404 1317 2444 1323
rect 2484 1317 2716 1323
rect 2724 1317 2764 1323
rect 2845 1323 2851 1337
rect 2868 1337 2908 1343
rect 2964 1337 2972 1343
rect 3076 1337 3180 1343
rect 3220 1337 3244 1343
rect 3460 1337 3484 1343
rect 3492 1337 3532 1343
rect 3604 1337 4044 1343
rect 4052 1337 4108 1343
rect 4180 1337 4220 1343
rect 4228 1337 4284 1343
rect 4436 1337 4764 1343
rect 4772 1337 4828 1343
rect 4980 1337 5052 1343
rect 5204 1337 5212 1343
rect 5252 1337 5436 1343
rect 5700 1337 5756 1343
rect 2845 1317 2876 1323
rect 2884 1317 2908 1323
rect 2973 1323 2979 1336
rect 2973 1317 3084 1323
rect 3188 1317 3228 1323
rect 3428 1317 3676 1323
rect 3892 1317 3948 1323
rect 4004 1317 4140 1323
rect 4148 1317 4156 1323
rect 4212 1317 4332 1323
rect 4436 1317 4556 1323
rect 4804 1317 4892 1323
rect 4900 1317 5004 1323
rect 5028 1317 5100 1323
rect 5316 1317 5580 1323
rect 5588 1317 5628 1323
rect 5645 1317 5660 1323
rect 5668 1317 5756 1323
rect 5876 1317 5964 1323
rect 5972 1317 6012 1323
rect 36 1297 108 1303
rect 276 1297 332 1303
rect 404 1297 460 1303
rect 468 1297 700 1303
rect 708 1297 780 1303
rect 820 1297 844 1303
rect 900 1297 940 1303
rect 964 1297 1004 1303
rect 1028 1297 1052 1303
rect 1060 1297 1244 1303
rect 1396 1297 1500 1303
rect 1508 1297 1532 1303
rect 1620 1297 1676 1303
rect 1748 1297 1804 1303
rect 2052 1297 2140 1303
rect 2164 1297 2236 1303
rect 2596 1297 2620 1303
rect 2740 1297 2780 1303
rect 2820 1297 2892 1303
rect 3028 1297 3212 1303
rect 3252 1297 3340 1303
rect 3757 1303 3763 1316
rect 3476 1297 3763 1303
rect 4036 1297 4252 1303
rect 4500 1297 4636 1303
rect 4772 1297 5084 1303
rect 5092 1297 5164 1303
rect 5348 1297 5420 1303
rect 5604 1297 5644 1303
rect 5812 1297 5900 1303
rect 6020 1297 6044 1303
rect 148 1277 172 1283
rect 292 1277 348 1283
rect 388 1277 444 1283
rect 884 1277 1180 1283
rect 1188 1277 1324 1283
rect 1556 1277 1644 1283
rect 1716 1277 1772 1283
rect 1972 1277 2236 1283
rect 2244 1277 2316 1283
rect 2420 1277 3500 1283
rect 3524 1277 3644 1283
rect 3716 1277 3820 1283
rect 3828 1277 3852 1283
rect 3860 1277 3900 1283
rect 4180 1277 4188 1283
rect 4324 1277 4460 1283
rect 4468 1277 4524 1283
rect 4532 1277 4716 1283
rect 5508 1277 5564 1283
rect 5572 1277 5612 1283
rect 180 1257 364 1263
rect 740 1257 1132 1263
rect 1396 1257 1612 1263
rect 1636 1257 1836 1263
rect 1876 1257 1996 1263
rect 2004 1257 2012 1263
rect 2036 1257 2524 1263
rect 2532 1257 2572 1263
rect 2628 1257 2748 1263
rect 2772 1257 3276 1263
rect 3300 1257 3340 1263
rect 3348 1257 3468 1263
rect 3501 1263 3507 1276
rect 3501 1257 4252 1263
rect 4260 1257 4300 1263
rect 4372 1257 4396 1263
rect 4484 1257 4844 1263
rect 4852 1257 5052 1263
rect 5364 1257 6012 1263
rect 308 1237 492 1243
rect 692 1237 924 1243
rect 1348 1237 1596 1243
rect 1940 1237 2204 1243
rect 2260 1237 2268 1243
rect 2308 1237 2796 1243
rect 2852 1237 2940 1243
rect 3172 1237 3660 1243
rect 3668 1237 3788 1243
rect 3908 1237 4364 1243
rect 4452 1237 5244 1243
rect 5252 1237 5292 1243
rect 532 1217 988 1223
rect 1092 1217 1388 1223
rect 2084 1217 2092 1223
rect 2148 1217 2396 1223
rect 2516 1217 2700 1223
rect 3380 1217 3532 1223
rect 3549 1217 3868 1223
rect 1560 1214 1608 1216
rect 1560 1206 1564 1214
rect 1574 1206 1580 1214
rect 1588 1206 1594 1214
rect 1604 1206 1608 1214
rect 1560 1204 1608 1206
rect 356 1197 396 1203
rect 692 1197 908 1203
rect 916 1197 1132 1203
rect 1300 1197 1324 1203
rect 1748 1197 1932 1203
rect 1940 1197 2188 1203
rect 2228 1197 2428 1203
rect 2500 1197 2812 1203
rect 2836 1197 3292 1203
rect 3549 1203 3555 1217
rect 3876 1217 3916 1223
rect 4180 1217 4204 1223
rect 4340 1217 4380 1223
rect 4632 1214 4680 1216
rect 4632 1206 4636 1214
rect 4646 1206 4652 1214
rect 4660 1206 4666 1214
rect 4676 1206 4680 1214
rect 4632 1204 4680 1206
rect 3332 1197 3555 1203
rect 3572 1197 3580 1203
rect 3604 1197 3628 1203
rect 3652 1197 3740 1203
rect 3764 1197 4028 1203
rect 4212 1197 4428 1203
rect -19 1177 -13 1183
rect 724 1177 764 1183
rect 804 1177 876 1183
rect 980 1177 1260 1183
rect 1460 1177 1555 1183
rect 628 1157 700 1163
rect 740 1157 860 1163
rect 1012 1157 1068 1163
rect 1412 1157 1436 1163
rect 1444 1157 1516 1163
rect 1549 1163 1555 1177
rect 1572 1177 1644 1183
rect 1652 1177 1756 1183
rect 1828 1177 1932 1183
rect 1956 1177 2172 1183
rect 2356 1177 2604 1183
rect 2708 1177 3084 1183
rect 3092 1177 3228 1183
rect 3236 1177 3308 1183
rect 3508 1177 3516 1183
rect 3572 1177 3596 1183
rect 3764 1177 3900 1183
rect 3924 1177 4012 1183
rect 4372 1177 4860 1183
rect 5156 1177 5244 1183
rect 1549 1157 1820 1163
rect 2349 1163 2355 1176
rect 1844 1157 2355 1163
rect 2404 1157 2620 1163
rect 2644 1157 2668 1163
rect 2676 1157 2860 1163
rect 2884 1157 3020 1163
rect 3060 1157 3196 1163
rect 3220 1157 3276 1163
rect 3405 1157 3564 1163
rect 3405 1144 3411 1157
rect 3572 1157 3612 1163
rect 3636 1157 3756 1163
rect 3933 1157 3996 1163
rect 548 1137 1116 1143
rect 1124 1137 1180 1143
rect 1204 1137 1228 1143
rect 1476 1137 1500 1143
rect 1508 1137 1596 1143
rect 1604 1137 1900 1143
rect 1940 1137 1948 1143
rect 2004 1137 2076 1143
rect 2084 1137 2124 1143
rect 2148 1137 2252 1143
rect 2356 1137 2444 1143
rect 2580 1137 2739 1143
rect 116 1117 188 1123
rect 212 1117 268 1123
rect 324 1117 348 1123
rect 356 1117 572 1123
rect 724 1117 812 1123
rect 820 1117 1068 1123
rect 1364 1117 1468 1123
rect 1476 1117 1708 1123
rect 1732 1117 1996 1123
rect 2020 1117 2092 1123
rect 2100 1117 2140 1123
rect 2164 1117 2220 1123
rect 2260 1117 2332 1123
rect 2436 1117 2444 1123
rect 2596 1117 2652 1123
rect 2733 1123 2739 1137
rect 2772 1137 2908 1143
rect 2932 1137 3244 1143
rect 3252 1137 3340 1143
rect 3364 1137 3404 1143
rect 3540 1137 3548 1143
rect 3588 1137 3692 1143
rect 3933 1143 3939 1157
rect 4404 1157 4940 1163
rect 4948 1157 4988 1163
rect 5188 1157 5692 1163
rect 3748 1137 3939 1143
rect 3956 1137 4076 1143
rect 4356 1137 5260 1143
rect 5268 1137 5340 1143
rect 5460 1137 5596 1143
rect 6285 1137 6291 1143
rect 2733 1117 2780 1123
rect 2788 1117 2892 1123
rect 2932 1117 2972 1123
rect 3028 1117 3100 1123
rect 3108 1117 3212 1123
rect 3268 1117 3308 1123
rect 3332 1117 3468 1123
rect 3540 1117 3596 1123
rect 3668 1117 3724 1123
rect 3780 1117 4188 1123
rect 4388 1117 4492 1123
rect 4500 1117 4636 1123
rect 4724 1117 4908 1123
rect 4916 1117 4956 1123
rect 5140 1117 5228 1123
rect 5732 1117 5916 1123
rect 100 1097 140 1103
rect 148 1097 156 1103
rect 164 1097 220 1103
rect 532 1097 588 1103
rect 596 1097 636 1103
rect 660 1097 844 1103
rect 852 1097 1052 1103
rect 1284 1097 1308 1103
rect 1428 1097 1452 1103
rect 1524 1097 1612 1103
rect 1645 1097 1676 1103
rect 116 1077 204 1083
rect 452 1077 508 1083
rect 580 1077 652 1083
rect 676 1077 812 1083
rect 820 1077 908 1083
rect 916 1077 956 1083
rect 980 1077 1164 1083
rect 1645 1083 1651 1097
rect 1684 1097 1740 1103
rect 1780 1097 1868 1103
rect 1892 1097 2508 1103
rect 2628 1097 2684 1103
rect 2740 1097 2796 1103
rect 2820 1097 2892 1103
rect 2916 1097 2988 1103
rect 3044 1097 3644 1103
rect 3652 1097 3708 1103
rect 3828 1097 3836 1103
rect 3908 1097 3916 1103
rect 3988 1097 4108 1103
rect 4260 1097 4412 1103
rect 4468 1097 4556 1103
rect 4564 1097 4780 1103
rect 4788 1097 4844 1103
rect 5044 1097 5052 1103
rect 5236 1097 5276 1103
rect 5284 1097 5372 1103
rect 5716 1097 5740 1103
rect 5796 1097 6108 1103
rect 1380 1077 1651 1083
rect 1668 1077 1724 1083
rect 1972 1077 2012 1083
rect 2132 1077 2140 1083
rect 2180 1077 2300 1083
rect 2356 1077 2380 1083
rect 2436 1077 2572 1083
rect 2580 1077 3180 1083
rect 3220 1077 3260 1083
rect 3300 1077 3324 1083
rect 3364 1077 3884 1083
rect 3892 1077 3980 1083
rect 3988 1077 4220 1083
rect 4292 1077 4547 1083
rect 84 1057 156 1063
rect 196 1057 412 1063
rect 756 1057 860 1063
rect 868 1057 988 1063
rect 1060 1057 1244 1063
rect 1492 1057 1708 1063
rect 1732 1057 1836 1063
rect 1908 1057 2348 1063
rect 2548 1057 3308 1063
rect 3332 1057 3372 1063
rect 3396 1057 3932 1063
rect 3940 1057 3948 1063
rect 4004 1057 4060 1063
rect 4084 1057 4252 1063
rect 4276 1057 4300 1063
rect 4541 1063 4547 1077
rect 4564 1077 4588 1083
rect 4836 1077 4892 1083
rect 4932 1077 5004 1083
rect 5268 1077 5324 1083
rect 5412 1077 5516 1083
rect 5524 1077 5580 1083
rect 5988 1077 6076 1083
rect 4541 1057 4732 1063
rect 4980 1057 5132 1063
rect 5284 1057 5660 1063
rect 5668 1057 5852 1063
rect 532 1037 668 1043
rect 676 1037 940 1043
rect 1044 1037 1116 1043
rect 1124 1037 1260 1043
rect 1709 1043 1715 1056
rect 1709 1037 1804 1043
rect 1956 1037 2172 1043
rect 2388 1037 2444 1043
rect 2484 1037 2956 1043
rect 2964 1037 3036 1043
rect 3044 1037 3068 1043
rect 3085 1037 3420 1043
rect 900 1017 972 1023
rect 980 1017 1020 1023
rect 1524 1017 1820 1023
rect 1828 1017 1852 1023
rect 2045 1017 2252 1023
rect 548 997 620 1003
rect 628 997 908 1003
rect 1028 997 1212 1003
rect 2045 1003 2051 1017
rect 2276 1017 2524 1023
rect 2740 1017 2764 1023
rect 3085 1023 3091 1037
rect 3444 1037 3500 1043
rect 3997 1043 4003 1056
rect 3556 1037 4003 1043
rect 4308 1037 4476 1043
rect 4484 1037 4748 1043
rect 4756 1037 4860 1043
rect 4996 1037 5196 1043
rect 5300 1037 5356 1043
rect 5364 1037 5404 1043
rect 5524 1037 5548 1043
rect 6052 1037 6204 1043
rect 2916 1017 3091 1023
rect 3437 1023 3443 1036
rect 3188 1017 3443 1023
rect 3492 1017 3564 1023
rect 3588 1017 3836 1023
rect 3860 1017 3884 1023
rect 4372 1017 4412 1023
rect 5140 1017 5244 1023
rect 5252 1017 5484 1023
rect 5556 1017 5628 1023
rect 5636 1017 5676 1023
rect 6196 1017 6236 1023
rect 3112 1014 3160 1016
rect 3112 1006 3116 1014
rect 3126 1006 3132 1014
rect 3140 1006 3146 1014
rect 3156 1006 3160 1014
rect 3112 1004 3160 1006
rect 1316 997 2051 1003
rect 2068 997 2236 1003
rect 2516 997 2556 1003
rect 2564 997 2588 1003
rect 3028 997 3084 1003
rect 3252 997 3260 1003
rect 3284 997 3443 1003
rect 132 977 332 983
rect 772 977 796 983
rect 852 977 1036 983
rect 1076 977 1148 983
rect 1412 977 1500 983
rect 1508 977 1708 983
rect 1716 977 1980 983
rect 2340 977 2412 983
rect 2420 977 2540 983
rect 2628 977 2860 983
rect 2868 977 3388 983
rect 3437 983 3443 997
rect 3460 997 4156 1003
rect 4564 997 4604 1003
rect 5044 997 5132 1003
rect 5140 997 5436 1003
rect 5492 997 5708 1003
rect 3437 977 3772 983
rect 3796 977 3820 983
rect 3844 977 3868 983
rect 3892 977 4012 983
rect 4036 977 4044 983
rect 4068 977 4444 983
rect 4548 977 4588 983
rect 4884 977 4908 983
rect 5060 977 5084 983
rect 5092 977 5116 983
rect 5188 977 5292 983
rect 5316 977 5404 983
rect 6036 977 6092 983
rect 6100 977 6156 983
rect -19 957 -13 963
rect 100 957 140 963
rect 212 957 243 963
rect 237 944 243 957
rect 276 957 284 963
rect 340 957 380 963
rect 436 957 492 963
rect 500 957 700 963
rect 740 957 812 963
rect 1076 957 1308 963
rect 1780 957 1820 963
rect 1828 957 1836 963
rect 1972 957 2028 963
rect 2084 957 2828 963
rect 2996 957 3036 963
rect 3044 957 3116 963
rect 3380 957 3436 963
rect 3444 957 3660 963
rect 3700 957 3852 963
rect 3860 957 3948 963
rect 3956 957 4092 963
rect 4180 957 4220 963
rect 4404 957 4428 963
rect 4468 957 4524 963
rect 4532 957 4700 963
rect 4708 957 4748 963
rect 4804 957 5020 963
rect 5028 957 5116 963
rect 5124 957 5148 963
rect 5652 957 5708 963
rect 52 937 108 943
rect 196 937 220 943
rect 244 937 348 943
rect 708 937 748 943
rect 788 937 1356 943
rect 1844 937 2092 943
rect 2292 937 2636 943
rect 2644 937 2668 943
rect 2676 937 3452 943
rect 3572 937 3708 943
rect 3732 937 3804 943
rect 3876 937 3916 943
rect 3924 937 3980 943
rect 3997 937 4044 943
rect 3997 924 4003 937
rect 4340 937 4380 943
rect 4388 937 4396 943
rect 4436 937 4476 943
rect 4532 937 4556 943
rect 4580 937 4844 943
rect 4852 937 4892 943
rect 4900 937 4956 943
rect 4980 937 5052 943
rect 5140 937 5148 943
rect 5204 937 5244 943
rect 5972 937 5996 943
rect 6244 937 6291 943
rect -19 917 -13 923
rect 84 917 332 923
rect 420 917 476 923
rect 484 917 636 923
rect 660 917 1084 923
rect 1156 917 1196 923
rect 1396 917 1420 923
rect 1892 917 1948 923
rect 2036 917 2156 923
rect 2228 917 2268 923
rect 2308 917 2316 923
rect 2420 917 2460 923
rect 2484 917 2604 923
rect 2612 917 2860 923
rect 2868 917 3180 923
rect 3236 917 3276 923
rect 3300 917 3404 923
rect 3524 917 3660 923
rect 3668 917 3788 923
rect 3940 917 3996 923
rect 4036 917 4172 923
rect 4692 917 4732 923
rect 4916 917 5004 923
rect 5076 917 5228 923
rect 5236 917 5340 923
rect 5396 917 5452 923
rect 5460 917 5500 923
rect 5588 917 5628 923
rect 5636 917 5676 923
rect 5748 917 5852 923
rect 6164 917 6188 923
rect 132 897 140 903
rect 148 897 332 903
rect 452 897 620 903
rect 1076 897 1100 903
rect 1140 897 1228 903
rect 1236 897 1260 903
rect 1332 897 1340 903
rect 1556 897 1660 903
rect 1668 897 1724 903
rect 1732 897 1788 903
rect 1844 897 1948 903
rect 1956 897 1996 903
rect 2212 897 2380 903
rect 2404 897 2524 903
rect 2596 897 2652 903
rect 2660 897 2860 903
rect 2900 897 2908 903
rect 2916 897 3436 903
rect 3604 897 3644 903
rect 3684 897 3804 903
rect 3812 897 3900 903
rect 4244 897 4348 903
rect 4468 897 4508 903
rect 4804 897 4860 903
rect 5005 903 5011 916
rect 5005 897 5100 903
rect 5220 897 5356 903
rect 5364 897 5532 903
rect 5636 897 5788 903
rect 5988 897 6092 903
rect 6148 897 6291 903
rect 36 877 76 883
rect 260 877 396 883
rect 564 877 604 883
rect 916 877 988 883
rect 996 877 1020 883
rect 1092 877 1116 883
rect 1124 877 1164 883
rect 1348 877 1372 883
rect 1396 877 1628 883
rect 1636 877 1740 883
rect 1748 877 1804 883
rect 1940 877 2188 883
rect 2340 877 2396 883
rect 2404 877 2492 883
rect 2548 877 2588 883
rect 2660 877 2796 883
rect 2932 877 2940 883
rect 2948 877 3036 883
rect 3060 877 3212 883
rect 3268 877 3724 883
rect 3748 877 3772 883
rect 3924 877 3980 883
rect 4740 877 4924 883
rect 5108 877 5180 883
rect 5396 877 5612 883
rect 5620 877 5660 883
rect 6100 877 6204 883
rect 676 857 1388 863
rect 1460 857 1484 863
rect 1620 857 1660 863
rect 1700 857 2044 863
rect 2052 857 2108 863
rect 2196 857 2684 863
rect 2692 857 2707 863
rect 2756 857 2780 863
rect 2932 857 3500 863
rect 3940 857 5468 863
rect 5476 857 5548 863
rect 628 837 684 843
rect 1332 837 1516 843
rect 1524 837 1564 843
rect 1572 837 1692 843
rect 1876 837 1948 843
rect 1972 837 2108 843
rect 2116 837 2172 843
rect 2180 837 2444 843
rect 2580 837 3020 843
rect 3460 837 5196 843
rect 5492 837 6060 843
rect 1108 817 1180 823
rect 2196 817 2364 823
rect 2708 817 2956 823
rect 2996 817 3052 823
rect 3092 817 3388 823
rect 3396 817 3404 823
rect 3812 817 4460 823
rect 5332 817 6156 823
rect 1560 814 1608 816
rect 1560 806 1564 814
rect 1574 806 1580 814
rect 1588 806 1594 814
rect 1604 806 1608 814
rect 1560 804 1608 806
rect 4632 814 4680 816
rect 4632 806 4636 814
rect 4646 806 4652 814
rect 4660 806 4666 814
rect 4676 806 4680 814
rect 4632 804 4680 806
rect 932 797 1100 803
rect 1108 797 1148 803
rect 1812 797 2012 803
rect 2036 797 2348 803
rect 2740 797 2748 803
rect 2804 797 3212 803
rect 4180 797 4204 803
rect 5364 797 5516 803
rect 244 777 300 783
rect 308 777 332 783
rect 500 777 588 783
rect 1028 777 1116 783
rect 1140 777 1228 783
rect 1428 777 1548 783
rect 1892 777 2156 783
rect 2388 777 2460 783
rect 2772 777 3308 783
rect 3316 777 3340 783
rect 3924 777 4332 783
rect 5924 777 5996 783
rect 324 757 652 763
rect 948 757 972 763
rect 1316 757 1756 763
rect 1876 757 2204 763
rect 2212 757 2348 763
rect 2436 757 2668 763
rect 2724 757 2796 763
rect 3044 757 3388 763
rect 3844 757 3900 763
rect 4820 757 4972 763
rect 6285 757 6291 763
rect 324 737 364 743
rect 372 737 412 743
rect 436 737 460 743
rect 500 737 540 743
rect 836 737 1036 743
rect 1300 737 1372 743
rect 1380 737 1468 743
rect 1476 737 1564 743
rect 1828 737 1884 743
rect 2100 737 2140 743
rect 2260 737 2444 743
rect 2500 737 2540 743
rect 2708 737 2764 743
rect 2852 737 3196 743
rect 3684 737 3708 743
rect 3732 737 3916 743
rect 3924 737 3964 743
rect 3988 737 4012 743
rect 4564 737 4700 743
rect 4756 737 4780 743
rect 4980 737 5292 743
rect 5300 737 5324 743
rect 5348 737 5468 743
rect 5476 737 5532 743
rect 5540 737 5580 743
rect 5780 737 5884 743
rect 5972 737 6188 743
rect 68 717 252 723
rect 388 717 684 723
rect 948 717 1068 723
rect 1172 717 1260 723
rect 1428 717 1820 723
rect 1860 717 2060 723
rect 2244 717 2364 723
rect 2372 717 2412 723
rect 2445 723 2451 736
rect 2445 717 2508 723
rect 2532 717 2700 723
rect 2708 717 2780 723
rect 2788 717 3356 723
rect 3412 717 3724 723
rect 3748 717 3788 723
rect 3828 717 4252 723
rect 4260 717 4300 723
rect 4452 717 4476 723
rect 4580 717 4668 723
rect 4852 717 5004 723
rect 5044 717 5084 723
rect 5172 717 5356 723
rect 5716 717 5916 723
rect 6228 717 6236 723
rect 84 697 172 703
rect 212 697 236 703
rect 292 697 348 703
rect 436 697 524 703
rect 580 697 620 703
rect 788 697 828 703
rect 1236 697 1452 703
rect 1460 697 1548 703
rect 1780 697 1980 703
rect 1988 697 2188 703
rect 2196 697 2220 703
rect 2228 697 2284 703
rect 2340 697 2796 703
rect 2804 697 2876 703
rect 2884 697 2924 703
rect 2964 697 3052 703
rect 3172 697 3292 703
rect 3300 697 3356 703
rect 3476 697 3532 703
rect 3540 697 3548 703
rect 3572 697 3644 703
rect 3668 697 3724 703
rect 3732 697 3772 703
rect 3780 697 3820 703
rect 3924 697 3948 703
rect 3956 697 3980 703
rect 4004 697 4156 703
rect 4372 697 4444 703
rect 4532 697 4556 703
rect 4612 697 4684 703
rect 4740 697 4796 703
rect 4804 697 4908 703
rect 5060 697 5212 703
rect 5300 697 5436 703
rect 5460 697 5500 703
rect 5668 697 5820 703
rect 6180 697 6291 703
rect 100 677 204 683
rect 228 677 444 683
rect 452 677 508 683
rect 772 677 812 683
rect 820 677 844 683
rect 932 677 988 683
rect 1076 677 1164 683
rect 1284 677 1340 683
rect 1748 677 1836 683
rect 1844 677 1900 683
rect 2116 677 2172 683
rect 2372 677 2812 683
rect 2820 677 2844 683
rect 2852 677 2908 683
rect 2980 677 3020 683
rect 3268 677 3596 683
rect 3620 677 4012 683
rect 4036 677 4044 683
rect 4148 677 4172 683
rect 4340 677 4396 683
rect 4548 677 4748 683
rect 4804 677 5260 683
rect 5268 677 5340 683
rect 5460 677 5548 683
rect 276 657 364 663
rect 404 657 588 663
rect 644 657 780 663
rect 1220 657 1292 663
rect 1396 657 1516 663
rect 2164 657 2332 663
rect 2612 657 2668 663
rect 2836 657 2972 663
rect 3076 657 3260 663
rect 3460 657 3516 663
rect 3588 657 3660 663
rect 3668 657 3804 663
rect 3812 657 3852 663
rect 4196 657 4540 663
rect 4596 657 4732 663
rect 4740 657 4876 663
rect 4884 657 4956 663
rect 5076 657 5228 663
rect 5236 657 5260 663
rect 5268 657 5404 663
rect 6180 657 6220 663
rect 6285 657 6291 663
rect 68 637 652 643
rect 669 637 924 643
rect 116 617 220 623
rect 669 623 675 637
rect 932 637 1004 643
rect 1220 637 1484 643
rect 1581 637 1948 643
rect 468 617 675 623
rect 804 617 1308 623
rect 1581 623 1587 637
rect 1956 637 2028 643
rect 2468 637 2508 643
rect 2532 637 2652 643
rect 2820 637 3276 643
rect 3284 637 3388 643
rect 3508 637 3532 643
rect 3588 637 3932 643
rect 4100 637 4380 643
rect 4404 637 5052 643
rect 5076 637 5100 643
rect 5124 637 5324 643
rect 5876 637 5964 643
rect 6132 637 6220 643
rect 1364 617 1587 623
rect 1604 617 1996 623
rect 2004 617 2140 623
rect 2148 617 2316 623
rect 2324 617 2380 623
rect 2692 617 2988 623
rect 3188 617 3276 623
rect 3284 617 3404 623
rect 3716 617 4524 623
rect 4548 617 4716 623
rect 4724 617 4796 623
rect 4980 617 5196 623
rect 5220 617 5340 623
rect 5908 617 5948 623
rect 3112 614 3160 616
rect 3112 606 3116 614
rect 3126 606 3132 614
rect 3140 606 3146 614
rect 3156 606 3160 614
rect 3112 604 3160 606
rect 260 597 524 603
rect 628 597 684 603
rect 836 597 1004 603
rect 1012 597 1068 603
rect 1364 597 1916 603
rect 2356 597 2508 603
rect 2676 597 2796 603
rect 2804 597 2892 603
rect 3956 597 4956 603
rect 5508 597 5804 603
rect 5812 597 5852 603
rect 100 577 140 583
rect 212 577 291 583
rect 100 557 268 563
rect 285 563 291 577
rect 340 577 604 583
rect 612 577 684 583
rect 692 577 716 583
rect 740 577 764 583
rect 788 577 1116 583
rect 1460 577 1612 583
rect 1684 577 1964 583
rect 1972 577 2012 583
rect 2260 577 2732 583
rect 2772 577 3148 583
rect 3165 577 3468 583
rect 285 557 460 563
rect 516 557 572 563
rect 580 557 636 563
rect 708 557 892 563
rect 980 557 1228 563
rect 1348 557 1420 563
rect 1540 557 2076 563
rect 2084 557 2092 563
rect 2404 557 2428 563
rect 2452 557 2508 563
rect 2548 557 2556 563
rect 2564 557 2604 563
rect 3165 563 3171 577
rect 3796 577 4044 583
rect 4052 577 4108 583
rect 4180 577 4236 583
rect 4276 577 4476 583
rect 4484 577 4556 583
rect 4564 577 4764 583
rect 4788 577 5116 583
rect 5124 577 5164 583
rect 5172 577 5212 583
rect 5396 577 5692 583
rect 5940 577 5964 583
rect 2852 557 3171 563
rect 3181 557 3244 563
rect 3181 544 3187 557
rect 3284 557 3420 563
rect 3508 557 3612 563
rect 3732 557 3836 563
rect 3844 557 3916 563
rect 3940 557 3980 563
rect 4292 557 4332 563
rect 4420 557 4460 563
rect 4628 557 5043 563
rect 116 537 380 543
rect 388 537 428 543
rect 644 537 700 543
rect 740 537 1132 543
rect 1140 537 1228 543
rect 1236 537 1292 543
rect 1316 537 1356 543
rect 1444 537 1772 543
rect 1780 537 2172 543
rect 2180 537 2268 543
rect 2532 537 2572 543
rect 2612 537 2780 543
rect 2788 537 2860 543
rect 2884 537 2940 543
rect 3012 537 3036 543
rect 3124 537 3180 543
rect 3252 537 3708 543
rect 3716 537 3820 543
rect 3876 537 3964 543
rect 4020 537 4076 543
rect 4132 537 4188 543
rect 4548 537 4636 543
rect 4772 537 4812 543
rect 4852 537 4972 543
rect 5037 543 5043 557
rect 5076 557 5484 563
rect 5492 557 5532 563
rect 5037 537 5132 543
rect 5204 537 5356 543
rect 5588 537 5836 543
rect 5844 537 5916 543
rect 276 517 316 523
rect 580 517 748 523
rect 900 517 956 523
rect 1124 517 1164 523
rect 1332 517 1484 523
rect 1508 517 1548 523
rect 1620 517 1676 523
rect 1844 517 1916 523
rect 2228 517 2396 523
rect 2516 517 2556 523
rect 3028 517 3068 523
rect 3076 517 3292 523
rect 3300 517 4204 523
rect 4212 517 4300 523
rect 4333 517 4364 523
rect 196 497 236 503
rect 285 497 332 503
rect 285 484 291 497
rect 397 497 492 503
rect 148 477 284 483
rect 397 483 403 497
rect 500 497 540 503
rect 564 497 652 503
rect 660 497 844 503
rect 1172 497 1692 503
rect 1700 497 1740 503
rect 1748 497 1788 503
rect 2164 497 2220 503
rect 2244 497 2284 503
rect 2532 497 3164 503
rect 3172 497 3212 503
rect 3284 497 3292 503
rect 3380 497 3468 503
rect 3476 497 3516 503
rect 4333 503 4339 517
rect 4372 517 4444 523
rect 4468 517 4508 523
rect 4532 517 4956 523
rect 5428 517 5500 523
rect 5588 517 5644 523
rect 5700 517 5740 523
rect 6164 517 6220 523
rect 3812 497 4339 503
rect 4356 497 4492 503
rect 4500 497 4588 503
rect 4596 497 4748 503
rect 4756 497 4860 503
rect 4980 497 5068 503
rect 5140 497 5180 503
rect 5396 497 5596 503
rect 5604 497 5628 503
rect 6180 497 6188 503
rect 6212 497 6291 503
rect 308 477 403 483
rect 420 477 476 483
rect 484 477 524 483
rect 692 477 716 483
rect 740 477 780 483
rect 1012 477 1660 483
rect 1668 477 1724 483
rect 1732 477 1772 483
rect 1892 477 1932 483
rect 1940 477 1980 483
rect 2036 477 2268 483
rect 2276 477 2380 483
rect 2724 477 2764 483
rect 2772 477 2956 483
rect 3172 477 3868 483
rect 3876 477 3900 483
rect 3908 477 3948 483
rect 4196 477 4332 483
rect 4484 477 5020 483
rect 5028 477 5468 483
rect 5476 477 5516 483
rect 5620 477 5772 483
rect 244 457 860 463
rect 996 457 1052 463
rect 1076 457 1340 463
rect 1380 457 1420 463
rect 1428 457 1628 463
rect 1636 457 1708 463
rect 1716 457 1756 463
rect 1764 457 1820 463
rect 1940 457 2620 463
rect 2628 457 2732 463
rect 2900 457 3260 463
rect 3268 457 3308 463
rect 3476 457 3852 463
rect 3892 457 4156 463
rect 5076 457 5100 463
rect 5428 457 6236 463
rect 84 437 124 443
rect 452 437 908 443
rect 1076 437 1388 443
rect 1412 437 1452 443
rect 1476 437 1852 443
rect 1860 437 1900 443
rect 2308 437 2812 443
rect 2948 437 3692 443
rect 4004 437 4380 443
rect 4388 437 4428 443
rect 4468 437 5084 443
rect 5092 437 5148 443
rect 5156 437 5308 443
rect 5332 437 5580 443
rect 5588 437 5708 443
rect -19 417 -13 423
rect 132 417 396 423
rect 500 417 828 423
rect 836 417 1116 423
rect 1124 417 1276 423
rect 1812 417 2540 423
rect 3684 417 4220 423
rect 4228 417 4252 423
rect 4372 417 4524 423
rect 4548 417 4572 423
rect 5108 417 5564 423
rect 5572 417 5676 423
rect 1560 414 1608 416
rect 1560 406 1564 414
rect 1574 406 1580 414
rect 1588 406 1594 414
rect 1604 406 1608 414
rect 1560 404 1608 406
rect 4632 414 4680 416
rect 4632 406 4636 414
rect 4646 406 4652 414
rect 4660 406 4666 414
rect 4676 406 4680 414
rect 4632 404 4680 406
rect 308 397 348 403
rect 356 397 396 403
rect 404 397 524 403
rect 548 397 684 403
rect 708 397 844 403
rect 932 397 1036 403
rect 1140 397 1500 403
rect 1652 397 1836 403
rect 2356 397 3004 403
rect 3700 397 3884 403
rect 3908 397 4012 403
rect 4036 397 4236 403
rect 4756 397 5244 403
rect 5364 397 5420 403
rect 5428 397 5612 403
rect 5908 397 5932 403
rect -19 377 -13 383
rect 52 377 92 383
rect 468 377 764 383
rect 772 377 1020 383
rect 1028 377 1244 383
rect 1700 377 2076 383
rect 2132 377 2444 383
rect 3364 377 3916 383
rect 3940 377 3980 383
rect 3988 377 4140 383
rect 276 357 460 363
rect 564 357 764 363
rect 788 357 1084 363
rect 1204 357 1372 363
rect 1492 357 1612 363
rect 1620 357 1676 363
rect 1892 357 1948 363
rect 2596 357 3788 363
rect 3796 357 3836 363
rect 4052 357 4124 363
rect 5252 357 5436 363
rect 5636 357 5740 363
rect 6212 357 6291 363
rect 260 337 492 343
rect 500 337 588 343
rect 596 337 812 343
rect 893 337 988 343
rect 52 317 140 323
rect 148 317 204 323
rect 484 317 572 323
rect 580 317 636 323
rect 660 317 732 323
rect 893 323 899 337
rect 1028 337 1068 343
rect 1092 337 1116 343
rect 1124 337 1180 343
rect 1268 337 1308 343
rect 1332 337 1388 343
rect 1524 337 1628 343
rect 1844 337 2236 343
rect 2804 337 2844 343
rect 2852 337 2908 343
rect 2916 337 3484 343
rect 3540 337 3660 343
rect 3956 337 4364 343
rect 4372 337 4476 343
rect 4916 337 4956 343
rect 5076 337 5260 343
rect 5341 337 5404 343
rect 5341 324 5347 337
rect 5588 337 5644 343
rect 5828 337 5916 343
rect 5924 337 6012 343
rect 772 317 899 323
rect 916 317 988 323
rect 1012 317 1212 323
rect 1220 317 1324 323
rect 1332 317 1340 323
rect 1748 317 2060 323
rect 2260 317 2428 323
rect 2436 317 2476 323
rect 2500 317 2636 323
rect 2724 317 2764 323
rect 2772 317 2812 323
rect 2836 317 2860 323
rect 3076 317 3212 323
rect 3332 317 3372 323
rect 3380 317 3420 323
rect 3437 317 3580 323
rect 68 297 124 303
rect 164 297 220 303
rect 324 297 364 303
rect 372 297 444 303
rect 516 297 556 303
rect 564 297 620 303
rect 692 297 716 303
rect 724 297 956 303
rect 980 297 1132 303
rect 1140 297 1196 303
rect 1252 297 1324 303
rect 1380 297 1436 303
rect 1444 297 1484 303
rect 1572 297 1788 303
rect 1828 297 1900 303
rect 2468 297 2556 303
rect 2660 297 2796 303
rect 2820 297 2892 303
rect 3437 303 3443 317
rect 3972 317 3980 323
rect 4004 317 4028 323
rect 4116 317 4140 323
rect 4324 317 4348 323
rect 4436 317 4556 323
rect 4564 317 4572 323
rect 4612 317 4780 323
rect 5140 317 5164 323
rect 5188 317 5340 323
rect 5396 317 5404 323
rect 5460 317 5516 323
rect 5556 317 6220 323
rect 6260 317 6291 323
rect 3396 297 3443 303
rect 3460 297 3500 303
rect 3668 297 3692 303
rect 3876 297 4620 303
rect 4628 297 4908 303
rect 4916 297 4940 303
rect 5044 297 5148 303
rect 5156 297 5228 303
rect 5332 297 5612 303
rect 5620 297 5756 303
rect 5828 297 5836 303
rect 5924 297 5996 303
rect 52 277 92 283
rect 212 277 252 283
rect 388 277 412 283
rect 420 277 556 283
rect 756 277 780 283
rect 868 277 1068 283
rect 1108 277 1244 283
rect 1284 277 1308 283
rect 1332 277 1724 283
rect 1860 277 2076 283
rect 2196 277 2284 283
rect 2292 277 2364 283
rect 2436 277 2604 283
rect 2612 277 2652 283
rect 2932 277 3148 283
rect 3236 277 3340 283
rect 3492 277 3708 283
rect 3956 277 3996 283
rect 4020 277 4028 283
rect 4100 277 4268 283
rect 4884 277 4924 283
rect 5012 277 5036 283
rect 5044 277 5068 283
rect 5076 277 5084 283
rect 5220 277 5500 283
rect 5508 277 5532 283
rect 5556 277 5580 283
rect 5668 277 5900 283
rect 5908 277 5964 283
rect 196 257 236 263
rect 372 257 652 263
rect 660 257 876 263
rect 884 257 1052 263
rect 1124 257 1452 263
rect 1460 257 1692 263
rect 1732 257 1932 263
rect 2164 257 2188 263
rect 2244 257 2316 263
rect 2324 257 2332 263
rect 2644 257 2748 263
rect 3524 257 3756 263
rect 3764 257 3804 263
rect 4020 257 4300 263
rect 4308 257 4444 263
rect 4452 257 4524 263
rect 4996 257 5052 263
rect 5533 263 5539 276
rect 5533 257 5660 263
rect 5668 257 5676 263
rect 5892 257 5932 263
rect 6004 257 6108 263
rect 356 237 540 243
rect 612 237 796 243
rect 820 237 924 243
rect 1028 237 1260 243
rect 1284 237 1356 243
rect 1396 237 1715 243
rect 180 217 236 223
rect 436 217 908 223
rect 916 217 972 223
rect 1012 217 1148 223
rect 1156 217 1228 223
rect 1268 217 1500 223
rect 1508 217 1596 223
rect 1709 223 1715 237
rect 1732 237 1852 243
rect 2452 237 2764 243
rect 2996 237 3036 243
rect 3044 237 3180 243
rect 3300 237 4076 243
rect 4148 237 4252 243
rect 4484 237 4636 243
rect 4820 237 4972 243
rect 4980 237 5356 243
rect 5444 237 5916 243
rect 1709 217 1788 223
rect 1796 217 1820 223
rect 1860 217 2108 223
rect 2420 217 2828 223
rect 3780 217 4588 223
rect 5412 217 5740 223
rect 3112 214 3160 216
rect 3112 206 3116 214
rect 3126 206 3132 214
rect 3140 206 3146 214
rect 3156 206 3160 214
rect 3112 204 3160 206
rect 148 197 412 203
rect 468 197 668 203
rect 868 197 1420 203
rect 1492 197 1564 203
rect 1748 197 2140 203
rect 2772 197 3084 203
rect 3540 197 3596 203
rect 3620 197 3900 203
rect 4020 197 4108 203
rect 4868 197 5132 203
rect 5556 197 5804 203
rect 5812 197 5868 203
rect 228 177 524 183
rect 532 177 588 183
rect 701 177 1164 183
rect 84 157 284 163
rect 701 163 707 177
rect 1501 177 1836 183
rect 1501 164 1507 177
rect 2484 177 4876 183
rect 4932 177 4988 183
rect 4996 177 5100 183
rect 5140 177 5308 183
rect 5316 177 5468 183
rect 5476 177 5676 183
rect 6132 177 6156 183
rect 548 157 707 163
rect 724 157 796 163
rect 820 157 988 163
rect 1012 157 1148 163
rect 1300 157 1372 163
rect 1444 157 1500 163
rect 1860 157 1916 163
rect 1924 157 1948 163
rect 1988 157 2028 163
rect 2052 157 2076 163
rect 2340 157 2380 163
rect 2388 157 2675 163
rect 196 137 364 143
rect 388 137 508 143
rect 516 137 556 143
rect 644 137 732 143
rect 740 137 812 143
rect 861 137 1228 143
rect 861 124 867 137
rect 1316 137 1340 143
rect 1412 137 1436 143
rect 1540 137 1628 143
rect 1924 137 2188 143
rect 2612 137 2652 143
rect 2669 143 2675 157
rect 2756 157 2812 163
rect 2900 157 2924 163
rect 3204 157 3308 163
rect 3508 157 3644 163
rect 3796 157 3868 163
rect 4148 157 4316 163
rect 4372 157 4428 163
rect 4852 157 4892 163
rect 4964 157 5148 163
rect 5204 157 5260 163
rect 5492 157 5644 163
rect 5908 157 5932 163
rect 6036 157 6220 163
rect 2669 137 3052 143
rect 3124 137 3452 143
rect 3652 137 3692 143
rect 3700 137 3788 143
rect 3860 137 4044 143
rect 4260 137 4300 143
rect 4308 137 4364 143
rect 4388 137 4460 143
rect 4532 137 4620 143
rect 4788 137 5996 143
rect 6068 137 6172 143
rect 84 117 188 123
rect 260 117 316 123
rect 324 117 396 123
rect 452 117 492 123
rect 660 117 748 123
rect 788 117 860 123
rect 948 117 1244 123
rect 1252 117 1516 123
rect 1892 117 2012 123
rect 2036 117 2044 123
rect 2196 117 2236 123
rect 2244 117 2348 123
rect 2532 117 2620 123
rect 2676 117 2700 123
rect 2724 117 2796 123
rect 2804 117 2908 123
rect 3076 117 3212 123
rect 3316 117 3340 123
rect 3460 117 3548 123
rect 3556 117 3660 123
rect 3748 117 3836 123
rect 3844 117 3932 123
rect 4756 117 4828 123
rect 4900 117 5004 123
rect 5076 117 5228 123
rect 5348 117 5420 123
rect 5444 117 5468 123
rect 5620 117 5708 123
rect 5780 117 5804 123
rect 5940 117 5987 123
rect 52 97 284 103
rect 292 97 332 103
rect 372 97 508 103
rect 516 97 604 103
rect 692 97 716 103
rect 740 97 764 103
rect 772 97 1100 103
rect 1364 97 1388 103
rect 1460 97 1484 103
rect 1956 97 1964 103
rect 1972 97 1996 103
rect 2621 103 2627 116
rect 2621 97 2764 103
rect 2788 97 2876 103
rect 2980 97 3052 103
rect 3188 97 3260 103
rect 3716 97 3788 103
rect 4292 97 4428 103
rect 4980 97 5084 103
rect 5316 97 5340 103
rect 5348 97 5420 103
rect 5572 97 5628 103
rect 5636 97 5644 103
rect 5876 97 5964 103
rect 5981 103 5987 117
rect 6004 117 6172 123
rect 5981 97 6028 103
rect 628 77 876 83
rect 884 77 908 83
rect 916 77 956 83
rect 1076 77 1116 83
rect 5380 77 5548 83
rect 5556 77 5596 83
rect 5620 77 5820 83
rect 292 57 844 63
rect 1069 63 1075 76
rect 932 57 1075 63
rect 2708 57 2780 63
rect 3444 57 3564 63
rect -19 37 -13 43
rect 3540 37 3564 43
rect 3860 37 4124 43
rect 4180 37 4252 43
rect 6285 37 6291 43
rect 2324 17 2332 23
rect 2516 17 2604 23
rect 3508 17 3532 23
rect 4820 17 4844 23
rect 5924 17 5964 23
rect 6164 17 6172 23
rect 1560 14 1608 16
rect 1560 6 1564 14
rect 1574 6 1580 14
rect 1588 6 1594 14
rect 1604 6 1608 14
rect 1560 4 1608 6
rect 4632 14 4680 16
rect 4632 6 4636 14
rect 4646 6 4652 14
rect 4660 6 4666 14
rect 4676 6 4680 14
rect 4632 4 4680 6
<< m4contact >>
rect 3116 5806 3118 5814
rect 3118 5806 3124 5814
rect 3132 5806 3140 5814
rect 3148 5806 3154 5814
rect 3154 5806 3156 5814
rect 1068 5796 1076 5804
rect 1132 5796 1140 5804
rect 3052 5796 3060 5804
rect 1964 5756 1972 5764
rect 588 5736 596 5744
rect 1068 5736 1076 5744
rect 5900 5736 5908 5744
rect 204 5716 212 5724
rect 908 5716 916 5724
rect 2028 5716 2036 5724
rect 2252 5696 2260 5704
rect 1452 5676 1460 5684
rect 6028 5676 6036 5684
rect 1132 5636 1140 5644
rect 5228 5636 5236 5644
rect 1564 5606 1566 5614
rect 1566 5606 1572 5614
rect 1580 5606 1588 5614
rect 1596 5606 1602 5614
rect 1602 5606 1604 5614
rect 4636 5606 4638 5614
rect 4638 5606 4644 5614
rect 4652 5606 4660 5614
rect 4668 5606 4674 5614
rect 4674 5606 4676 5614
rect 3724 5596 3732 5604
rect 5548 5576 5556 5584
rect 460 5536 468 5544
rect 2796 5536 2804 5544
rect 5196 5536 5204 5544
rect 6252 5536 6260 5544
rect 1260 5516 1268 5524
rect 1356 5516 1364 5524
rect 1452 5516 1460 5524
rect 5452 5516 5460 5524
rect 6092 5496 6100 5504
rect 12 5476 20 5484
rect 2380 5476 2388 5484
rect 2700 5476 2708 5484
rect 3948 5476 3956 5484
rect 6156 5476 6164 5484
rect 204 5456 212 5464
rect 620 5456 628 5464
rect 1516 5456 1524 5464
rect 5388 5456 5396 5464
rect 396 5436 404 5444
rect 588 5436 596 5444
rect 1036 5436 1044 5444
rect 1420 5416 1428 5424
rect 3756 5436 3764 5444
rect 3116 5406 3118 5414
rect 3118 5406 3124 5414
rect 3132 5406 3140 5414
rect 3148 5406 3154 5414
rect 3154 5406 3156 5414
rect 972 5396 980 5404
rect 5644 5396 5652 5404
rect 5900 5396 5908 5404
rect 460 5376 468 5384
rect 1260 5376 1268 5384
rect 3564 5376 3572 5384
rect 12 5336 20 5344
rect 2284 5356 2292 5364
rect 908 5336 916 5344
rect 1420 5336 1428 5344
rect 3500 5336 3508 5344
rect 4588 5336 4596 5344
rect 5836 5336 5844 5344
rect 6220 5336 6228 5344
rect 3692 5316 3700 5324
rect 396 5296 404 5304
rect 5932 5316 5940 5324
rect 6124 5316 6132 5324
rect 6220 5296 6228 5304
rect 620 5276 628 5284
rect 1068 5276 1076 5284
rect 2700 5276 2708 5284
rect 2796 5276 2804 5284
rect 3692 5276 3700 5284
rect 1356 5256 1364 5264
rect 5132 5256 5140 5264
rect 2284 5236 2292 5244
rect 4044 5236 4052 5244
rect 6188 5236 6196 5244
rect 5580 5216 5588 5224
rect 6252 5216 6260 5224
rect 1564 5206 1566 5214
rect 1566 5206 1572 5214
rect 1580 5206 1588 5214
rect 1596 5206 1602 5214
rect 1602 5206 1604 5214
rect 4636 5206 4638 5214
rect 4638 5206 4644 5214
rect 4652 5206 4660 5214
rect 4668 5206 4674 5214
rect 4674 5206 4676 5214
rect 140 5176 148 5184
rect 3564 5176 3572 5184
rect 3948 5176 3956 5184
rect 4364 5156 4372 5164
rect 5740 5136 5748 5144
rect 3468 5116 3476 5124
rect 5964 5116 5972 5124
rect 908 5076 916 5084
rect 5196 5096 5204 5104
rect 6252 5096 6260 5104
rect 1420 5076 1428 5084
rect 3580 5076 3588 5084
rect 4588 5076 4596 5084
rect 76 5056 84 5064
rect 2636 5056 2644 5064
rect 3884 5056 3892 5064
rect 6060 5056 6068 5064
rect 6220 5056 6228 5064
rect 3500 5036 3508 5044
rect 3852 5036 3860 5044
rect 5772 5036 5780 5044
rect 2508 5016 2516 5024
rect 3116 5006 3118 5014
rect 3118 5006 3124 5014
rect 3132 5006 3140 5014
rect 3148 5006 3154 5014
rect 3154 5006 3156 5014
rect 1260 4996 1268 5004
rect 1676 4996 1684 5004
rect 1804 4996 1812 5004
rect 5964 4976 5972 4984
rect 6124 4976 6132 4984
rect 6220 4976 6228 4984
rect 844 4936 852 4944
rect 972 4936 980 4944
rect 1036 4936 1044 4944
rect 3084 4936 3092 4944
rect 3404 4936 3412 4944
rect 3852 4936 3860 4944
rect 4460 4936 4468 4944
rect 4908 4936 4916 4944
rect 6028 4936 6036 4944
rect 2508 4916 2516 4924
rect 4044 4916 4052 4924
rect 4204 4916 4212 4924
rect 5260 4916 5268 4924
rect 5964 4916 5972 4924
rect 3052 4896 3060 4904
rect 3372 4896 3380 4904
rect 4908 4896 4916 4904
rect 3532 4876 3540 4884
rect 5132 4876 5140 4884
rect 6028 4876 6036 4884
rect 6220 4876 6228 4884
rect 556 4836 564 4844
rect 1564 4806 1566 4814
rect 1566 4806 1572 4814
rect 1580 4806 1588 4814
rect 1596 4806 1602 4814
rect 1602 4806 1604 4814
rect 4636 4806 4638 4814
rect 4638 4806 4644 4814
rect 4652 4806 4660 4814
rect 4668 4806 4674 4814
rect 4674 4806 4676 4814
rect 1196 4796 1204 4804
rect 5292 4796 5300 4804
rect 812 4756 820 4764
rect 972 4756 980 4764
rect 1388 4756 1396 4764
rect 2380 4756 2388 4764
rect 3052 4756 3060 4764
rect 5004 4756 5012 4764
rect 4396 4736 4404 4744
rect 5932 4736 5940 4744
rect 2732 4716 2740 4724
rect 4044 4716 4052 4724
rect 3436 4696 3444 4704
rect 3852 4696 3860 4704
rect 5868 4696 5876 4704
rect 6092 4696 6100 4704
rect 6220 4696 6228 4704
rect 652 4676 660 4684
rect 2028 4676 2036 4684
rect 108 4656 116 4664
rect 908 4656 916 4664
rect 2636 4656 2644 4664
rect 3756 4656 3764 4664
rect 3820 4656 3828 4664
rect 5388 4656 5396 4664
rect 5900 4656 5908 4664
rect 6156 4656 6164 4664
rect 140 4636 148 4644
rect 204 4636 212 4644
rect 940 4636 948 4644
rect 1292 4636 1300 4644
rect 5516 4636 5524 4644
rect 3884 4616 3892 4624
rect 3116 4606 3118 4614
rect 3118 4606 3124 4614
rect 3132 4606 3140 4614
rect 3148 4606 3154 4614
rect 3154 4606 3156 4614
rect 4396 4596 4404 4604
rect 12 4576 20 4584
rect 1036 4576 1044 4584
rect 3756 4556 3764 4564
rect 12 4536 20 4544
rect 5132 4536 5140 4544
rect 76 4516 84 4524
rect 492 4516 500 4524
rect 5228 4536 5236 4544
rect 6124 4536 6132 4544
rect 6156 4536 6164 4544
rect 5260 4516 5268 4524
rect 5292 4516 5300 4524
rect 5644 4516 5652 4524
rect 652 4496 660 4504
rect 3084 4496 3092 4504
rect 3596 4496 3604 4504
rect 4588 4496 4596 4504
rect 4908 4496 4916 4504
rect 5388 4496 5396 4504
rect 44 4476 52 4484
rect 684 4476 692 4484
rect 2476 4476 2484 4484
rect 2732 4476 2740 4484
rect 3052 4476 3060 4484
rect 3276 4476 3284 4484
rect 3532 4476 3540 4484
rect 5932 4476 5940 4484
rect 2380 4456 2388 4464
rect 2892 4456 2900 4464
rect 3372 4456 3380 4464
rect 3436 4456 3444 4464
rect 4492 4456 4500 4464
rect 4204 4436 4212 4444
rect 4460 4436 4468 4444
rect 6028 4436 6036 4444
rect 6124 4436 6132 4444
rect 5708 4416 5716 4424
rect 1564 4406 1566 4414
rect 1566 4406 1572 4414
rect 1580 4406 1588 4414
rect 1596 4406 1602 4414
rect 1602 4406 1604 4414
rect 4636 4406 4638 4414
rect 4638 4406 4644 4414
rect 4652 4406 4660 4414
rect 4668 4406 4674 4414
rect 4674 4406 4676 4414
rect 3372 4376 3380 4384
rect 5740 4376 5748 4384
rect 1036 4356 1044 4364
rect 1644 4356 1652 4364
rect 3404 4356 3412 4364
rect 6028 4356 6036 4364
rect 44 4336 52 4344
rect 204 4336 212 4344
rect 2988 4336 2996 4344
rect 3436 4336 3444 4344
rect 5164 4336 5172 4344
rect 5580 4336 5588 4344
rect 5804 4336 5812 4344
rect 6092 4336 6100 4344
rect 5356 4316 5364 4324
rect 5740 4316 5748 4324
rect 460 4296 468 4304
rect 2220 4296 2228 4304
rect 2956 4296 2964 4304
rect 3276 4296 3284 4304
rect 5164 4296 5172 4304
rect 5644 4296 5652 4304
rect 172 4276 180 4284
rect 332 4276 340 4284
rect 588 4276 596 4284
rect 4460 4276 4468 4284
rect 684 4256 692 4264
rect 1100 4256 1108 4264
rect 2220 4256 2228 4264
rect 2668 4256 2676 4264
rect 3564 4256 3572 4264
rect 3628 4256 3636 4264
rect 5132 4256 5140 4264
rect 5292 4256 5300 4264
rect 5452 4276 5460 4284
rect 6124 4276 6132 4284
rect 5964 4256 5972 4264
rect 364 4236 372 4244
rect 556 4236 564 4244
rect 1196 4236 1204 4244
rect 4044 4236 4052 4244
rect 4588 4236 4596 4244
rect 5708 4236 5716 4244
rect 5740 4236 5748 4244
rect 6124 4236 6132 4244
rect 6252 4256 6260 4264
rect 3116 4206 3118 4214
rect 3118 4206 3124 4214
rect 3132 4206 3140 4214
rect 3148 4206 3154 4214
rect 3154 4206 3156 4214
rect 1132 4196 1140 4204
rect 4236 4196 4244 4204
rect 4748 4196 4756 4204
rect 5388 4196 5396 4204
rect 5452 4196 5460 4204
rect 5644 4176 5652 4184
rect 5964 4196 5972 4204
rect 1292 4156 1300 4164
rect 1356 4156 1364 4164
rect 2252 4156 2260 4164
rect 2380 4156 2388 4164
rect 3276 4156 3284 4164
rect 5356 4156 5364 4164
rect 524 4136 532 4144
rect 844 4136 852 4144
rect 1132 4116 1140 4124
rect 2252 4116 2260 4124
rect 5676 4136 5684 4144
rect 6092 4176 6100 4184
rect 3660 4116 3668 4124
rect 4876 4116 4884 4124
rect 364 4096 372 4104
rect 492 4096 500 4104
rect 844 4096 852 4104
rect 940 4096 948 4104
rect 1388 4096 1396 4104
rect 2668 4096 2676 4104
rect 2892 4096 2900 4104
rect 2956 4096 2964 4104
rect 3340 4096 3348 4104
rect 4268 4096 4276 4104
rect 4332 4096 4340 4104
rect 4492 4096 4500 4104
rect 5164 4116 5172 4124
rect 5452 4116 5460 4124
rect 5804 4136 5812 4144
rect 6124 4136 6132 4144
rect 6252 4156 6260 4164
rect 3372 4076 3380 4084
rect 4460 4076 4468 4084
rect 5644 4096 5652 4104
rect 5420 4076 5428 4084
rect 5484 4076 5492 4084
rect 5676 4076 5684 4084
rect 6092 4096 6100 4104
rect 6124 4096 6132 4104
rect 6252 4096 6260 4104
rect 588 4056 596 4064
rect 2604 4056 2612 4064
rect 2988 4056 2996 4064
rect 3596 4056 3604 4064
rect 4748 4056 4756 4064
rect 5164 4056 5172 4064
rect 5996 4056 6004 4064
rect 3468 4036 3476 4044
rect 3756 4036 3764 4044
rect 4876 4036 4884 4044
rect 5388 4036 5396 4044
rect 5516 4036 5524 4044
rect 5452 4016 5460 4024
rect 1564 4006 1566 4014
rect 1566 4006 1572 4014
rect 1580 4006 1588 4014
rect 1596 4006 1602 4014
rect 1602 4006 1604 4014
rect 4636 4006 4638 4014
rect 4638 4006 4644 4014
rect 4652 4006 4660 4014
rect 4668 4006 4674 4014
rect 4674 4006 4676 4014
rect 172 3996 180 4004
rect 4748 3996 4756 4004
rect 2028 3976 2036 3984
rect 12 3956 20 3964
rect 5356 3956 5364 3964
rect 6252 3936 6260 3944
rect 3852 3916 3860 3924
rect 4588 3916 4596 3924
rect 5708 3916 5716 3924
rect 6124 3916 6132 3924
rect 3436 3896 3444 3904
rect 5260 3896 5268 3904
rect 5324 3896 5332 3904
rect 12 3876 20 3884
rect 652 3876 660 3884
rect 1036 3876 1044 3884
rect 1164 3876 1172 3884
rect 1324 3876 1332 3884
rect 2636 3876 2644 3884
rect 4236 3876 4244 3884
rect 4268 3876 4276 3884
rect 4332 3876 4340 3884
rect 5292 3876 5300 3884
rect 6124 3876 6132 3884
rect 684 3856 692 3864
rect 1100 3856 1108 3864
rect 3212 3856 3220 3864
rect 1132 3836 1140 3844
rect 1836 3836 1844 3844
rect 2604 3836 2612 3844
rect 3180 3836 3188 3844
rect 3276 3836 3284 3844
rect 3564 3856 3572 3864
rect 5612 3856 5620 3864
rect 4012 3836 4020 3844
rect 5276 3836 5284 3844
rect 332 3816 340 3824
rect 620 3816 628 3824
rect 1324 3816 1332 3824
rect 2252 3816 2260 3824
rect 3500 3816 3508 3824
rect 3116 3806 3118 3814
rect 3118 3806 3124 3814
rect 3132 3806 3140 3814
rect 3148 3806 3154 3814
rect 3154 3806 3156 3814
rect 3084 3796 3092 3804
rect 3852 3796 3860 3804
rect 5132 3796 5140 3804
rect 5932 3796 5940 3804
rect 844 3776 852 3784
rect 1420 3776 1428 3784
rect 3308 3776 3316 3784
rect 3564 3776 3572 3784
rect 3596 3776 3604 3784
rect 5292 3776 5300 3784
rect 5644 3776 5652 3784
rect 2636 3756 2644 3764
rect 3340 3756 3348 3764
rect 6252 3776 6260 3784
rect 172 3736 180 3744
rect 1292 3736 1300 3744
rect 2604 3736 2612 3744
rect 3660 3736 3668 3744
rect 5612 3736 5620 3744
rect 5804 3736 5812 3744
rect 6028 3736 6036 3744
rect 6252 3736 6260 3744
rect 108 3716 116 3724
rect 844 3716 852 3724
rect 1356 3716 1364 3724
rect 1452 3716 1460 3724
rect 3052 3716 3060 3724
rect 3596 3716 3604 3724
rect 5228 3716 5236 3724
rect 5516 3716 5524 3724
rect 492 3696 500 3704
rect 780 3696 788 3704
rect 876 3696 884 3704
rect 1132 3696 1140 3704
rect 1324 3696 1332 3704
rect 3084 3696 3092 3704
rect 5644 3696 5652 3704
rect 5900 3696 5908 3704
rect 5932 3696 5940 3704
rect 44 3676 52 3684
rect 268 3676 276 3684
rect 364 3676 372 3684
rect 1356 3676 1364 3684
rect 1388 3676 1396 3684
rect 3500 3676 3508 3684
rect 5996 3676 6004 3684
rect 1164 3656 1172 3664
rect 1228 3656 1236 3664
rect 1644 3656 1652 3664
rect 4204 3656 4212 3664
rect 6124 3676 6132 3684
rect 556 3636 564 3644
rect 716 3636 724 3644
rect 940 3636 948 3644
rect 1836 3636 1844 3644
rect 2860 3636 2868 3644
rect 4460 3636 4468 3644
rect 1260 3616 1268 3624
rect 2476 3616 2484 3624
rect 3340 3616 3348 3624
rect 1564 3606 1566 3614
rect 1566 3606 1572 3614
rect 1580 3606 1588 3614
rect 1596 3606 1602 3614
rect 1602 3606 1604 3614
rect 4636 3606 4638 3614
rect 4638 3606 4644 3614
rect 4652 3606 4660 3614
rect 4668 3606 4674 3614
rect 4674 3606 4676 3614
rect 492 3596 500 3604
rect 1804 3596 1812 3604
rect 2924 3596 2932 3604
rect 3276 3596 3284 3604
rect 6188 3616 6196 3624
rect 6252 3596 6260 3604
rect 2604 3576 2612 3584
rect 6060 3576 6068 3584
rect 460 3556 468 3564
rect 1356 3556 1364 3564
rect 2316 3556 2324 3564
rect 4140 3556 4148 3564
rect 2956 3536 2964 3544
rect 5932 3536 5940 3544
rect 6060 3536 6068 3544
rect 6124 3536 6132 3544
rect 1644 3516 1652 3524
rect 2252 3516 2260 3524
rect 3692 3516 3700 3524
rect 3724 3516 3732 3524
rect 4748 3516 4756 3524
rect 140 3496 148 3504
rect 1820 3476 1828 3484
rect 3532 3496 3540 3504
rect 5548 3496 5556 3504
rect 1964 3476 1972 3484
rect 3020 3476 3028 3484
rect 3404 3476 3412 3484
rect 3500 3476 3508 3484
rect 716 3436 724 3444
rect 1196 3436 1204 3444
rect 2892 3456 2900 3464
rect 4140 3456 4148 3464
rect 6252 3476 6260 3484
rect 2252 3436 2260 3444
rect 2668 3436 2676 3444
rect 2924 3436 2932 3444
rect 2956 3436 2964 3444
rect 5260 3436 5268 3444
rect 5292 3436 5300 3444
rect 940 3416 948 3424
rect 2604 3416 2612 3424
rect 5068 3416 5076 3424
rect 6124 3416 6132 3424
rect 3116 3406 3118 3414
rect 3118 3406 3124 3414
rect 3132 3406 3140 3414
rect 3148 3406 3154 3414
rect 3154 3406 3156 3414
rect 236 3396 244 3404
rect 748 3396 756 3404
rect 1484 3396 1492 3404
rect 2316 3396 2324 3404
rect 364 3376 372 3384
rect 1740 3376 1748 3384
rect 3756 3396 3764 3404
rect 5580 3396 5588 3404
rect 3436 3376 3444 3384
rect 3628 3376 3636 3384
rect 3692 3376 3700 3384
rect 5676 3376 5684 3384
rect 876 3356 884 3364
rect 1036 3356 1044 3364
rect 1868 3356 1876 3364
rect 2828 3356 2836 3364
rect 3052 3356 3060 3364
rect 3564 3356 3572 3364
rect 3660 3356 3668 3364
rect 6124 3356 6132 3364
rect 236 3336 244 3344
rect 588 3336 596 3344
rect 716 3336 724 3344
rect 908 3336 916 3344
rect 1292 3336 1300 3344
rect 300 3296 308 3304
rect 1004 3316 1012 3324
rect 1068 3316 1076 3324
rect 1100 3316 1108 3324
rect 1452 3316 1460 3324
rect 1228 3296 1236 3304
rect 1388 3296 1396 3304
rect 1484 3316 1492 3324
rect 4492 3336 4500 3344
rect 5068 3336 5076 3344
rect 3404 3316 3412 3324
rect 3532 3316 3540 3324
rect 4844 3316 4852 3324
rect 5516 3316 5524 3324
rect 5708 3316 5716 3324
rect 5900 3316 5908 3324
rect 5964 3316 5972 3324
rect 6188 3316 6196 3324
rect 3372 3296 3380 3304
rect 3852 3296 3860 3304
rect 4908 3296 4916 3304
rect 204 3276 212 3284
rect 620 3276 628 3284
rect 940 3276 948 3284
rect 1644 3276 1652 3284
rect 2828 3276 2836 3284
rect 5708 3276 5716 3284
rect 5740 3276 5748 3284
rect 1676 3256 1684 3264
rect 1964 3256 1972 3264
rect 524 3236 532 3244
rect 5484 3236 5492 3244
rect 748 3216 756 3224
rect 1292 3216 1300 3224
rect 3500 3216 3508 3224
rect 3756 3216 3764 3224
rect 6028 3216 6036 3224
rect 6156 3216 6164 3224
rect 1564 3206 1566 3214
rect 1566 3206 1572 3214
rect 1580 3206 1588 3214
rect 1596 3206 1602 3214
rect 1602 3206 1604 3214
rect 4636 3206 4638 3214
rect 4638 3206 4644 3214
rect 4652 3206 4660 3214
rect 4668 3206 4674 3214
rect 4674 3206 4676 3214
rect 1068 3196 1076 3204
rect 1132 3196 1140 3204
rect 1452 3196 1460 3204
rect 1932 3196 1940 3204
rect 3212 3196 3220 3204
rect 5964 3196 5972 3204
rect 6060 3196 6068 3204
rect 5164 3176 5172 3184
rect 268 3156 276 3164
rect 332 3156 340 3164
rect 780 3156 788 3164
rect 876 3156 884 3164
rect 1772 3156 1780 3164
rect 1996 3156 2004 3164
rect 3436 3156 3444 3164
rect 5996 3156 6004 3164
rect 3276 3136 3284 3144
rect 4204 3136 4212 3144
rect 5420 3136 5428 3144
rect 6060 3136 6068 3144
rect 1836 3116 1844 3124
rect 3020 3116 3028 3124
rect 3244 3116 3252 3124
rect 3340 3116 3348 3124
rect 5740 3116 5748 3124
rect 5996 3116 6004 3124
rect 6028 3116 6036 3124
rect 3788 3096 3796 3104
rect 5708 3096 5716 3104
rect 236 3076 244 3084
rect 524 3076 532 3084
rect 2860 3076 2868 3084
rect 3564 3076 3572 3084
rect 3756 3076 3764 3084
rect 4460 3076 4468 3084
rect 4492 3076 4500 3084
rect 5452 3076 5460 3084
rect 5836 3076 5844 3084
rect 140 3056 148 3064
rect 556 3056 564 3064
rect 620 3056 628 3064
rect 1004 3056 1012 3064
rect 1068 3056 1076 3064
rect 2892 3056 2900 3064
rect 3276 3056 3284 3064
rect 3596 3056 3604 3064
rect 3628 3056 3636 3064
rect 3788 3056 3796 3064
rect 4076 3056 4084 3064
rect 4588 3056 4596 3064
rect 5772 3056 5780 3064
rect 172 3036 180 3044
rect 876 3036 884 3044
rect 1452 3036 1460 3044
rect 2924 3036 2932 3044
rect 3212 3036 3220 3044
rect 3724 3036 3732 3044
rect 4012 3036 4020 3044
rect 5964 3036 5972 3044
rect 300 3016 308 3024
rect 2796 3016 2804 3024
rect 3756 3016 3764 3024
rect 5004 3016 5012 3024
rect 5164 3016 5172 3024
rect 5292 3016 5300 3024
rect 5388 3016 5396 3024
rect 5772 3016 5780 3024
rect 3116 3006 3118 3014
rect 3118 3006 3124 3014
rect 3132 3006 3140 3014
rect 3148 3006 3154 3014
rect 3154 3006 3156 3014
rect 332 2996 340 3004
rect 1164 2996 1172 3004
rect 108 2976 116 2984
rect 3916 2996 3924 3004
rect 4492 2976 4500 2984
rect 5932 2976 5940 2984
rect 492 2956 500 2964
rect 748 2956 756 2964
rect 1324 2956 1332 2964
rect 1836 2956 1844 2964
rect 2860 2956 2868 2964
rect 2956 2956 2964 2964
rect 4140 2956 4148 2964
rect 5100 2956 5108 2964
rect 5260 2956 5268 2964
rect 5324 2956 5332 2964
rect 5356 2956 5364 2964
rect 5516 2956 5524 2964
rect 5708 2956 5716 2964
rect 6092 2956 6100 2964
rect 524 2936 532 2944
rect 940 2936 948 2944
rect 1068 2936 1076 2944
rect 1516 2936 1524 2944
rect 3564 2936 3572 2944
rect 3756 2936 3764 2944
rect 5804 2936 5812 2944
rect 5964 2936 5972 2944
rect 108 2916 116 2924
rect 652 2916 660 2924
rect 1164 2916 1172 2924
rect 3372 2916 3380 2924
rect 3724 2916 3732 2924
rect 556 2896 564 2904
rect 2700 2896 2708 2904
rect 4204 2896 4212 2904
rect 4300 2896 4308 2904
rect 4332 2896 4340 2904
rect 5036 2916 5044 2924
rect 5260 2916 5268 2924
rect 5388 2916 5396 2924
rect 5580 2916 5588 2924
rect 5356 2896 5364 2904
rect 5644 2896 5652 2904
rect 5996 2916 6004 2924
rect 6060 2916 6068 2924
rect 6220 2916 6228 2924
rect 5932 2896 5940 2904
rect 620 2876 628 2884
rect 940 2876 948 2884
rect 3276 2876 3284 2884
rect 1036 2856 1044 2864
rect 3692 2856 3700 2864
rect 3756 2856 3764 2864
rect 4556 2876 4564 2884
rect 4972 2876 4980 2884
rect 3916 2856 3924 2864
rect 5548 2856 5556 2864
rect 5644 2856 5652 2864
rect 5740 2856 5748 2864
rect 5804 2856 5812 2864
rect 6124 2856 6132 2864
rect 6156 2856 6164 2864
rect 236 2836 244 2844
rect 1164 2836 1172 2844
rect 1420 2836 1428 2844
rect 1708 2836 1716 2844
rect 3372 2836 3380 2844
rect 76 2816 84 2824
rect 364 2816 372 2824
rect 460 2816 468 2824
rect 2796 2816 2804 2824
rect 3468 2816 3476 2824
rect 3500 2816 3508 2824
rect 3884 2816 3892 2824
rect 4172 2816 4180 2824
rect 5420 2816 5428 2824
rect 1564 2806 1566 2814
rect 1566 2806 1572 2814
rect 1580 2806 1588 2814
rect 1596 2806 1602 2814
rect 1602 2806 1604 2814
rect 4636 2806 4638 2814
rect 4638 2806 4644 2814
rect 4652 2806 4660 2814
rect 4668 2806 4674 2814
rect 4674 2806 4676 2814
rect 2764 2796 2772 2804
rect 2956 2796 2964 2804
rect 3084 2796 3092 2804
rect 1772 2776 1780 2784
rect 3372 2776 3380 2784
rect 428 2756 436 2764
rect 588 2756 596 2764
rect 1644 2756 1652 2764
rect 780 2736 788 2744
rect 972 2736 980 2744
rect 1388 2736 1396 2744
rect 1420 2736 1428 2744
rect 2828 2736 2836 2744
rect 4204 2756 4212 2764
rect 4716 2756 4724 2764
rect 5068 2756 5076 2764
rect 5100 2756 5108 2764
rect 5484 2756 5492 2764
rect 5996 2756 6004 2764
rect 140 2716 148 2724
rect 652 2716 660 2724
rect 812 2716 820 2724
rect 1228 2716 1236 2724
rect 1964 2716 1972 2724
rect 2860 2716 2868 2724
rect 3404 2736 3412 2744
rect 3628 2736 3636 2744
rect 5740 2736 5748 2744
rect 6124 2736 6132 2744
rect 3468 2716 3476 2724
rect 4044 2716 4052 2724
rect 1260 2696 1268 2704
rect 3628 2696 3636 2704
rect 3756 2696 3764 2704
rect 3916 2696 3924 2704
rect 4588 2696 4596 2704
rect 4780 2716 4788 2724
rect 5100 2716 5108 2724
rect 5132 2716 5140 2724
rect 5900 2716 5908 2724
rect 6060 2716 6068 2724
rect 6092 2716 6100 2724
rect 4812 2696 4820 2704
rect 5996 2696 6004 2704
rect 204 2676 212 2684
rect 716 2676 724 2684
rect 1100 2676 1108 2684
rect 1708 2676 1716 2684
rect 2060 2676 2068 2684
rect 2732 2676 2740 2684
rect 3212 2676 3220 2684
rect 3468 2676 3476 2684
rect 4172 2676 4180 2684
rect 6092 2676 6100 2684
rect 6124 2676 6132 2684
rect 1132 2656 1140 2664
rect 1932 2656 1940 2664
rect 2796 2656 2804 2664
rect 3500 2656 3508 2664
rect 428 2636 436 2644
rect 2732 2636 2740 2644
rect 2988 2636 2996 2644
rect 1004 2616 1012 2624
rect 3788 2656 3796 2664
rect 3884 2656 3892 2664
rect 4076 2656 4084 2664
rect 5452 2656 5460 2664
rect 5484 2656 5492 2664
rect 5932 2656 5940 2664
rect 3340 2616 3348 2624
rect 4300 2636 4308 2644
rect 4940 2636 4948 2644
rect 5612 2636 5620 2644
rect 5740 2636 5748 2644
rect 3788 2616 3796 2624
rect 4172 2616 4180 2624
rect 5132 2616 5140 2624
rect 5580 2616 5588 2624
rect 6188 2636 6196 2644
rect 5900 2616 5908 2624
rect 3116 2606 3118 2614
rect 3118 2606 3124 2614
rect 3132 2606 3140 2614
rect 3148 2606 3154 2614
rect 3154 2606 3156 2614
rect 940 2596 948 2604
rect 1164 2596 1172 2604
rect 1356 2596 1364 2604
rect 3596 2596 3604 2604
rect 524 2576 532 2584
rect 1196 2576 1204 2584
rect 1068 2556 1076 2564
rect 1228 2556 1236 2564
rect 3532 2576 3540 2584
rect 3692 2576 3700 2584
rect 4044 2576 4052 2584
rect 3180 2556 3188 2564
rect 5356 2556 5364 2564
rect 5996 2576 6004 2584
rect 6028 2556 6036 2564
rect 524 2536 532 2544
rect 780 2536 788 2544
rect 844 2536 852 2544
rect 1324 2536 1332 2544
rect 2508 2536 2516 2544
rect 140 2516 148 2524
rect 684 2496 692 2504
rect 1228 2496 1236 2504
rect 1516 2516 1524 2524
rect 2828 2516 2836 2524
rect 3372 2536 3380 2544
rect 3404 2536 3412 2544
rect 3628 2536 3636 2544
rect 4204 2536 4212 2544
rect 3308 2516 3316 2524
rect 4012 2516 4020 2524
rect 4332 2536 4340 2544
rect 5036 2536 5044 2544
rect 5228 2536 5236 2544
rect 5260 2536 5268 2544
rect 5676 2536 5684 2544
rect 4588 2516 4596 2524
rect 5388 2516 5396 2524
rect 6124 2516 6132 2524
rect 6188 2516 6196 2524
rect 2924 2496 2932 2504
rect 2956 2496 2964 2504
rect 3788 2496 3796 2504
rect 3852 2496 3860 2504
rect 5132 2496 5140 2504
rect 5804 2496 5812 2504
rect 6156 2496 6164 2504
rect 364 2476 372 2484
rect 460 2476 468 2484
rect 492 2476 500 2484
rect 972 2476 980 2484
rect 1708 2476 1716 2484
rect 2860 2476 2868 2484
rect 3468 2476 3476 2484
rect 3532 2476 3540 2484
rect 4972 2476 4980 2484
rect 5964 2476 5972 2484
rect 1420 2456 1428 2464
rect 1740 2456 1748 2464
rect 3372 2456 3380 2464
rect 3916 2456 3924 2464
rect 4044 2456 4052 2464
rect 4076 2456 4084 2464
rect 108 2436 116 2444
rect 2636 2436 2644 2444
rect 4172 2436 4180 2444
rect 428 2416 436 2424
rect 1068 2416 1076 2424
rect 1996 2416 2004 2424
rect 2252 2416 2260 2424
rect 2604 2416 2612 2424
rect 2956 2416 2964 2424
rect 2988 2416 2996 2424
rect 3436 2416 3444 2424
rect 3756 2416 3764 2424
rect 3820 2416 3828 2424
rect 4556 2436 4564 2444
rect 4780 2436 4788 2444
rect 4876 2436 4884 2444
rect 6060 2436 6068 2444
rect 6092 2436 6100 2444
rect 6124 2436 6132 2444
rect 1564 2406 1566 2414
rect 1566 2406 1572 2414
rect 1580 2406 1588 2414
rect 1596 2406 1602 2414
rect 1602 2406 1604 2414
rect 4636 2406 4638 2414
rect 4638 2406 4644 2414
rect 4652 2406 4660 2414
rect 4668 2406 4674 2414
rect 4674 2406 4676 2414
rect 12 2396 20 2404
rect 396 2396 404 2404
rect 3052 2396 3060 2404
rect 3244 2396 3252 2404
rect 3340 2396 3348 2404
rect 3884 2396 3892 2404
rect 3948 2396 3956 2404
rect 6060 2396 6068 2404
rect 76 2376 84 2384
rect 108 2376 116 2384
rect 236 2356 244 2364
rect 364 2356 372 2364
rect 1388 2376 1396 2384
rect 2700 2376 2708 2384
rect 3820 2376 3828 2384
rect 4492 2376 4500 2384
rect 4972 2376 4980 2384
rect 5100 2376 5108 2384
rect 5260 2376 5268 2384
rect 5388 2376 5396 2384
rect 5580 2376 5588 2384
rect 5804 2376 5812 2384
rect 5900 2376 5908 2384
rect 1676 2356 1684 2364
rect 2508 2356 2516 2364
rect 3276 2356 3284 2364
rect 4172 2356 4180 2364
rect 5420 2356 5428 2364
rect 6028 2356 6036 2364
rect 6156 2356 6164 2364
rect 620 2336 628 2344
rect 2636 2336 2644 2344
rect 2668 2336 2676 2344
rect 3468 2336 3476 2344
rect 3916 2336 3924 2344
rect 4908 2336 4916 2344
rect 5100 2336 5108 2344
rect 5740 2336 5748 2344
rect 556 2316 564 2324
rect 588 2316 596 2324
rect 1132 2316 1140 2324
rect 1356 2316 1364 2324
rect 428 2296 436 2304
rect 748 2296 756 2304
rect 1516 2296 1524 2304
rect 2860 2296 2868 2304
rect 3020 2316 3028 2324
rect 3532 2316 3540 2324
rect 4396 2316 4404 2324
rect 5292 2316 5300 2324
rect 5356 2316 5364 2324
rect 5484 2316 5492 2324
rect 5900 2316 5908 2324
rect 5932 2316 5940 2324
rect 3180 2296 3188 2304
rect 3244 2296 3252 2304
rect 140 2276 148 2284
rect 1132 2276 1140 2284
rect 1420 2276 1428 2284
rect 2060 2276 2068 2284
rect 3020 2276 3028 2284
rect 3308 2276 3316 2284
rect 3340 2296 3348 2304
rect 3404 2296 3412 2304
rect 4492 2296 4500 2304
rect 4588 2296 4596 2304
rect 5804 2296 5812 2304
rect 5996 2296 6004 2304
rect 4556 2276 4564 2284
rect 4812 2276 4820 2284
rect 4940 2276 4948 2284
rect 5132 2276 5140 2284
rect 5420 2276 5428 2284
rect 5612 2276 5620 2284
rect 268 2256 276 2264
rect 300 2256 308 2264
rect 2604 2256 2612 2264
rect 332 2236 340 2244
rect 492 2236 500 2244
rect 1004 2236 1012 2244
rect 6156 2256 6164 2264
rect 5644 2236 5652 2244
rect 5900 2236 5908 2244
rect 6092 2236 6100 2244
rect 492 2196 500 2204
rect 2924 2216 2932 2224
rect 5964 2216 5972 2224
rect 6028 2216 6036 2224
rect 3116 2206 3118 2214
rect 3118 2206 3124 2214
rect 3132 2206 3140 2214
rect 3148 2206 3154 2214
rect 3154 2206 3156 2214
rect 2508 2196 2516 2204
rect 2892 2196 2900 2204
rect 3372 2196 3380 2204
rect 2252 2176 2260 2184
rect 3564 2176 3572 2184
rect 4428 2196 4436 2204
rect 3756 2176 3764 2184
rect 5740 2196 5748 2204
rect 6092 2196 6100 2204
rect 6156 2196 6164 2204
rect 5708 2176 5716 2184
rect 3052 2156 3060 2164
rect 3340 2156 3348 2164
rect 3468 2156 3476 2164
rect 5484 2156 5492 2164
rect 5612 2156 5620 2164
rect 2348 2136 2356 2144
rect 3020 2136 3028 2144
rect 3500 2136 3508 2144
rect 108 2096 116 2104
rect 748 2096 756 2104
rect 1644 2116 1652 2124
rect 2828 2116 2836 2124
rect 3244 2116 3252 2124
rect 2316 2096 2324 2104
rect 396 2076 404 2084
rect 876 2076 884 2084
rect 140 2056 148 2064
rect 2956 2076 2964 2084
rect 3404 2076 3412 2084
rect 5100 2136 5108 2144
rect 5996 2136 6004 2144
rect 4556 2116 4564 2124
rect 4844 2096 4852 2104
rect 6092 2116 6100 2124
rect 6124 2116 6132 2124
rect 1644 2056 1652 2064
rect 2476 2056 2484 2064
rect 2604 2056 2612 2064
rect 2860 2056 2868 2064
rect 3180 2056 3188 2064
rect 3372 2056 3380 2064
rect 3948 2076 3956 2084
rect 4108 2076 4116 2084
rect 5964 2096 5972 2104
rect 4044 2056 4052 2064
rect 4140 2056 4148 2064
rect 4716 2056 4724 2064
rect 4748 2056 4756 2064
rect 4972 2056 4980 2064
rect 5164 2056 5172 2064
rect 236 2036 244 2044
rect 1132 2036 1140 2044
rect 3020 2036 3028 2044
rect 76 2016 84 2024
rect 3180 2016 3188 2024
rect 4012 2016 4020 2024
rect 4396 2036 4404 2044
rect 4428 2036 4436 2044
rect 5132 2036 5140 2044
rect 6092 2036 6100 2044
rect 4748 2016 4756 2024
rect 5612 2016 5620 2024
rect 1564 2006 1566 2014
rect 1566 2006 1572 2014
rect 1580 2006 1588 2014
rect 1596 2006 1602 2014
rect 1602 2006 1604 2014
rect 4636 2006 4638 2014
rect 4638 2006 4644 2014
rect 4652 2006 4660 2014
rect 4668 2006 4674 2014
rect 4674 2006 4676 2014
rect 300 1996 308 2004
rect 588 1996 596 2004
rect 620 1996 628 2004
rect 1484 1996 1492 2004
rect 2412 1996 2420 2004
rect 3532 1996 3540 2004
rect 3820 1996 3828 2004
rect 4812 1996 4820 2004
rect 4844 1996 4852 2004
rect 5932 1996 5940 2004
rect 6028 1996 6036 2004
rect 556 1976 564 1984
rect 1644 1976 1652 1984
rect 3052 1976 3060 1984
rect 5068 1976 5076 1984
rect 6124 1976 6132 1984
rect 1164 1956 1172 1964
rect 2924 1956 2932 1964
rect 364 1936 372 1944
rect 492 1936 500 1944
rect 2060 1936 2068 1944
rect 908 1916 916 1924
rect 1164 1916 1172 1924
rect 2348 1936 2356 1944
rect 2444 1936 2452 1944
rect 2764 1936 2772 1944
rect 2124 1916 2132 1924
rect 3692 1936 3700 1944
rect 3948 1936 3956 1944
rect 5516 1936 5524 1944
rect 5708 1936 5716 1944
rect 4236 1916 4244 1924
rect 5644 1916 5652 1924
rect 6124 1916 6132 1924
rect 524 1896 532 1904
rect 844 1896 852 1904
rect 2348 1896 2356 1904
rect 4812 1896 4820 1904
rect 5932 1896 5940 1904
rect 6156 1896 6164 1904
rect 6220 1896 6228 1904
rect 12 1876 20 1884
rect 684 1876 692 1884
rect 716 1876 724 1884
rect 3276 1876 3284 1884
rect 3564 1876 3572 1884
rect 4108 1876 4116 1884
rect 492 1856 500 1864
rect 2348 1856 2356 1864
rect 812 1836 820 1844
rect 1484 1836 1492 1844
rect 2444 1856 2452 1864
rect 2956 1856 2964 1864
rect 3180 1856 3188 1864
rect 3596 1856 3604 1864
rect 2380 1836 2388 1844
rect 4524 1856 4532 1864
rect 4716 1856 4724 1864
rect 6028 1876 6036 1884
rect 6124 1876 6132 1884
rect 5900 1856 5908 1864
rect 6188 1856 6196 1864
rect 3788 1836 3796 1844
rect 5996 1836 6004 1844
rect 236 1816 244 1824
rect 268 1816 276 1824
rect 908 1816 916 1824
rect 1036 1816 1044 1824
rect 4012 1816 4020 1824
rect 3116 1806 3118 1814
rect 3118 1806 3124 1814
rect 3132 1806 3140 1814
rect 3148 1806 3154 1814
rect 3154 1806 3156 1814
rect 140 1776 148 1784
rect 652 1796 660 1804
rect 940 1796 948 1804
rect 2508 1796 2516 1804
rect 3084 1796 3092 1804
rect 3180 1796 3188 1804
rect 3884 1796 3892 1804
rect 4172 1796 4180 1804
rect 4716 1796 4724 1804
rect 5196 1796 5204 1804
rect 5804 1796 5812 1804
rect 5932 1796 5940 1804
rect 460 1776 468 1784
rect 1164 1776 1172 1784
rect 1388 1776 1396 1784
rect 1676 1776 1684 1784
rect 1932 1776 1940 1784
rect 2476 1776 2484 1784
rect 2796 1776 2804 1784
rect 3276 1776 3284 1784
rect 3308 1776 3316 1784
rect 3500 1776 3508 1784
rect 844 1736 852 1744
rect 908 1736 916 1744
rect 1260 1756 1268 1764
rect 2348 1756 2356 1764
rect 2604 1756 2612 1764
rect 3084 1756 3092 1764
rect 3692 1756 3700 1764
rect 3756 1756 3764 1764
rect 5036 1776 5044 1784
rect 4780 1756 4788 1764
rect 1068 1736 1076 1744
rect 1932 1736 1940 1744
rect 2060 1736 2068 1744
rect 332 1716 340 1724
rect 652 1716 660 1724
rect 684 1716 692 1724
rect 1132 1716 1140 1724
rect 1292 1716 1300 1724
rect 3020 1736 3028 1744
rect 3052 1736 3060 1744
rect 3180 1736 3188 1744
rect 3212 1736 3220 1744
rect 3660 1736 3668 1744
rect 5836 1736 5844 1744
rect 1868 1716 1876 1724
rect 3404 1716 3412 1724
rect 460 1696 468 1704
rect 524 1696 532 1704
rect 2604 1696 2612 1704
rect 3724 1696 3732 1704
rect 3916 1696 3924 1704
rect 4108 1696 4116 1704
rect 4140 1696 4148 1704
rect 4236 1696 4244 1704
rect 4876 1696 4884 1704
rect 5836 1696 5844 1704
rect 1100 1676 1108 1684
rect 5548 1676 5556 1684
rect 5868 1676 5876 1684
rect 6124 1676 6132 1684
rect 44 1656 52 1664
rect 1164 1656 1172 1664
rect 3020 1656 3028 1664
rect 3436 1656 3444 1664
rect 1516 1636 1524 1644
rect 1996 1636 2004 1644
rect 3756 1656 3764 1664
rect 4044 1636 4052 1644
rect 332 1616 340 1624
rect 492 1616 500 1624
rect 524 1616 532 1624
rect 652 1616 660 1624
rect 972 1616 980 1624
rect 1564 1606 1566 1614
rect 1566 1606 1572 1614
rect 1580 1606 1588 1614
rect 1596 1606 1602 1614
rect 1602 1606 1604 1614
rect 684 1596 692 1604
rect 5900 1616 5908 1624
rect 4636 1606 4638 1614
rect 4638 1606 4644 1614
rect 4652 1606 4660 1614
rect 4668 1606 4674 1614
rect 4674 1606 4676 1614
rect 3756 1596 3764 1604
rect 4108 1596 4116 1604
rect 4140 1596 4148 1604
rect 5260 1596 5268 1604
rect 844 1576 852 1584
rect 2444 1576 2452 1584
rect 3212 1576 3220 1584
rect 5900 1576 5908 1584
rect 2796 1556 2804 1564
rect 2988 1556 2996 1564
rect 3980 1556 3988 1564
rect 4812 1556 4820 1564
rect 5388 1556 5396 1564
rect 1228 1536 1236 1544
rect 2956 1536 2964 1544
rect 3852 1536 3860 1544
rect 716 1516 724 1524
rect 780 1516 788 1524
rect 812 1516 820 1524
rect 1036 1516 1044 1524
rect 2348 1516 2356 1524
rect 2604 1516 2612 1524
rect 524 1496 532 1504
rect 1196 1496 1204 1504
rect 1452 1496 1460 1504
rect 3276 1516 3284 1524
rect 3468 1516 3476 1524
rect 3884 1516 3892 1524
rect 5868 1516 5876 1524
rect 3180 1496 3188 1504
rect 3436 1496 3444 1504
rect 4780 1496 4788 1504
rect 5996 1496 6004 1504
rect 940 1476 948 1484
rect 1068 1476 1076 1484
rect 1228 1476 1236 1484
rect 2156 1476 2164 1484
rect 2668 1476 2676 1484
rect 3276 1476 3284 1484
rect 3564 1476 3572 1484
rect 4204 1476 4212 1484
rect 4460 1476 4468 1484
rect 5772 1476 5780 1484
rect 6156 1476 6164 1484
rect 972 1456 980 1464
rect 1292 1456 1300 1464
rect 2508 1456 2516 1464
rect 3180 1456 3188 1464
rect 6028 1456 6036 1464
rect 3788 1436 3796 1444
rect 588 1416 596 1424
rect 1836 1416 1844 1424
rect 2956 1416 2964 1424
rect 2988 1416 2996 1424
rect 3052 1416 3060 1424
rect 3276 1416 3284 1424
rect 3116 1406 3118 1414
rect 3118 1406 3124 1414
rect 3132 1406 3140 1414
rect 3148 1406 3154 1414
rect 3154 1406 3156 1414
rect 1004 1396 1012 1404
rect 2796 1396 2804 1404
rect 556 1376 564 1384
rect 620 1376 628 1384
rect 844 1376 852 1384
rect 972 1376 980 1384
rect 1196 1376 1204 1384
rect 3948 1416 3956 1424
rect 6060 1416 6068 1424
rect 3404 1376 3412 1384
rect 3532 1376 3540 1384
rect 3564 1376 3572 1384
rect 3692 1376 3700 1384
rect 4556 1376 4564 1384
rect 44 1356 52 1364
rect 108 1356 116 1364
rect 236 1356 244 1364
rect 1644 1356 1652 1364
rect 2092 1356 2100 1364
rect 780 1336 788 1344
rect 812 1336 820 1344
rect 1036 1336 1044 1344
rect 1452 1336 1460 1344
rect 588 1316 596 1324
rect 748 1316 756 1324
rect 972 1316 980 1324
rect 2668 1356 2676 1364
rect 3084 1356 3092 1364
rect 3788 1356 3796 1364
rect 5036 1356 5044 1364
rect 5644 1356 5652 1364
rect 2444 1316 2452 1324
rect 2956 1336 2964 1344
rect 3180 1336 3188 1344
rect 3212 1336 3220 1344
rect 3244 1336 3252 1344
rect 4044 1336 4052 1344
rect 4428 1336 4436 1344
rect 4972 1336 4980 1344
rect 5196 1336 5204 1344
rect 3692 1316 3700 1324
rect 3724 1316 3732 1324
rect 3756 1316 3764 1324
rect 4140 1316 4148 1324
rect 844 1296 852 1304
rect 1004 1296 1012 1304
rect 1388 1296 1396 1304
rect 2732 1296 2740 1304
rect 3020 1296 3028 1304
rect 3468 1296 3476 1304
rect 1644 1276 1652 1284
rect 1708 1276 1716 1284
rect 3660 1276 3668 1284
rect 4172 1276 4180 1284
rect 1996 1256 2004 1264
rect 2764 1256 2772 1264
rect 3340 1256 3348 1264
rect 4364 1256 4372 1264
rect 4396 1256 4404 1264
rect 4844 1256 4852 1264
rect 5356 1256 5364 1264
rect 1932 1236 1940 1244
rect 2252 1236 2260 1244
rect 524 1216 532 1224
rect 2092 1216 2100 1224
rect 2924 1216 2932 1224
rect 1564 1206 1566 1214
rect 1566 1206 1572 1214
rect 1580 1206 1588 1214
rect 1596 1206 1602 1214
rect 1602 1206 1604 1214
rect 1132 1196 1140 1204
rect 1292 1196 1300 1204
rect 4332 1216 4340 1224
rect 4636 1206 4638 1214
rect 4638 1206 4644 1214
rect 4652 1206 4660 1214
rect 4668 1206 4674 1214
rect 4674 1206 4676 1214
rect 3564 1196 3572 1204
rect 3628 1196 3636 1204
rect 4428 1196 4436 1204
rect 876 1176 884 1184
rect 940 1176 948 1184
rect 620 1156 628 1164
rect 1932 1176 1940 1184
rect 3500 1176 3508 1184
rect 3596 1176 3604 1184
rect 3212 1156 3220 1164
rect 3276 1156 3284 1164
rect 1196 1136 1204 1144
rect 1932 1136 1940 1144
rect 716 1116 724 1124
rect 1708 1116 1716 1124
rect 2444 1116 2452 1124
rect 3532 1136 3540 1144
rect 3948 1136 3956 1144
rect 140 1096 148 1104
rect 108 1076 116 1084
rect 812 1076 820 1084
rect 3820 1096 3828 1104
rect 3916 1096 3924 1104
rect 3980 1096 3988 1104
rect 5036 1096 5044 1104
rect 2124 1076 2132 1084
rect 2348 1076 2356 1084
rect 3884 1076 3892 1084
rect 76 1056 84 1064
rect 1484 1056 1492 1064
rect 1836 1056 1844 1064
rect 3308 1056 3316 1064
rect 3948 1056 3956 1064
rect 4556 1076 4564 1084
rect 5260 1076 5268 1084
rect 2476 1036 2484 1044
rect 428 996 436 1004
rect 2252 1016 2260 1024
rect 2764 1016 2772 1024
rect 5516 1036 5524 1044
rect 3468 1016 3476 1024
rect 6188 1016 6196 1024
rect 3116 1006 3118 1014
rect 3118 1006 3124 1014
rect 3132 1006 3140 1014
rect 3148 1006 3154 1014
rect 3154 1006 3156 1014
rect 2508 996 2516 1004
rect 2988 996 2996 1004
rect 3244 996 3252 1004
rect 1068 976 1076 984
rect 4556 996 4564 1004
rect 5132 996 5140 1004
rect 3788 976 3796 984
rect 3884 976 3892 984
rect 4012 976 4020 984
rect 4044 976 4052 984
rect 268 956 276 964
rect 332 956 340 964
rect 940 956 948 964
rect 2828 956 2836 964
rect 2988 956 2996 964
rect 3660 956 3668 964
rect 4172 956 4180 964
rect 2668 936 2676 944
rect 3724 936 3732 944
rect 3980 936 3988 944
rect 4396 936 4404 944
rect 4972 936 4980 944
rect 5132 936 5140 944
rect 2156 916 2164 924
rect 2316 916 2324 924
rect 2412 916 2420 924
rect 2604 916 2612 924
rect 3180 916 3188 924
rect 4172 916 4180 924
rect 6156 916 6164 924
rect 332 896 340 904
rect 1324 896 1332 904
rect 2380 896 2388 904
rect 2860 896 2868 904
rect 2892 896 2900 904
rect 3436 896 3444 904
rect 3596 896 3604 904
rect 2924 876 2932 884
rect 3212 876 3220 884
rect 3724 876 3732 884
rect 6092 876 6100 884
rect 1388 856 1396 864
rect 2444 836 2452 844
rect 3020 836 3028 844
rect 5484 836 5492 844
rect 6060 836 6068 844
rect 2956 816 2964 824
rect 2988 816 2996 824
rect 3052 816 3060 824
rect 4460 816 4468 824
rect 5324 816 5332 824
rect 6156 816 6164 824
rect 1564 806 1566 814
rect 1566 806 1572 814
rect 1580 806 1588 814
rect 1596 806 1602 814
rect 1602 806 1604 814
rect 4636 806 4638 814
rect 4638 806 4644 814
rect 4652 806 4660 814
rect 4668 806 4674 814
rect 4674 806 4676 814
rect 2348 796 2356 804
rect 2732 796 2740 804
rect 4172 796 4180 804
rect 4204 796 4212 804
rect 5356 796 5364 804
rect 3916 776 3924 784
rect 4332 776 4340 784
rect 3500 736 3508 744
rect 3980 736 3988 744
rect 5580 736 5588 744
rect 5964 736 5972 744
rect 1324 716 1332 724
rect 2700 716 2708 724
rect 3724 716 3732 724
rect 3788 716 3796 724
rect 3820 716 3828 724
rect 5036 716 5044 724
rect 5516 716 5524 724
rect 6220 716 6228 724
rect 236 696 244 704
rect 3532 696 3540 704
rect 4044 676 4052 684
rect 4748 676 4756 684
rect 268 656 276 664
rect 2412 656 2420 664
rect 2476 656 2484 664
rect 5260 656 5268 664
rect 460 616 468 624
rect 1484 636 1492 644
rect 5068 636 5076 644
rect 6124 636 6132 644
rect 2988 616 2996 624
rect 3276 616 3284 624
rect 4524 616 4532 624
rect 5900 616 5908 624
rect 3116 606 3118 614
rect 3118 606 3124 614
rect 3132 606 3140 614
rect 3148 606 3154 614
rect 3154 606 3156 614
rect 1356 596 1364 604
rect 2508 596 2516 604
rect 268 556 276 564
rect 1324 576 1332 584
rect 1452 576 1460 584
rect 3468 576 3476 584
rect 5388 576 5396 584
rect 5964 576 5972 584
rect 3980 556 3988 564
rect 428 536 436 544
rect 556 496 564 504
rect 652 496 660 504
rect 3276 496 3284 504
rect 4524 516 4532 524
rect 6156 516 6164 524
rect 6188 496 6196 504
rect 3468 456 3476 464
rect 5420 456 5428 464
rect 1452 436 1460 444
rect 1564 406 1566 414
rect 1566 406 1572 414
rect 1580 406 1588 414
rect 1596 406 1602 414
rect 1602 406 1604 414
rect 4636 406 4638 414
rect 4638 406 4644 414
rect 4652 406 4660 414
rect 4668 406 4674 414
rect 4674 406 4676 414
rect 524 396 532 404
rect 3884 396 3892 404
rect 4748 396 4756 404
rect 5900 396 5908 404
rect 5932 396 5940 404
rect 3916 376 3924 384
rect 460 356 468 364
rect 5580 336 5588 344
rect 1324 316 1332 324
rect 2828 316 2836 324
rect 2796 296 2804 304
rect 3980 316 3988 324
rect 4556 316 4564 324
rect 5388 316 5396 324
rect 5548 316 5556 324
rect 6252 316 6260 324
rect 5836 296 5844 304
rect 556 276 564 284
rect 1068 276 1076 284
rect 4012 276 4020 284
rect 5068 276 5076 284
rect 2156 256 2164 264
rect 2316 256 2324 264
rect 812 236 820 244
rect 1356 236 1364 244
rect 4076 236 4084 244
rect 5356 236 5364 244
rect 3116 206 3118 214
rect 3118 206 3124 214
rect 3132 206 3140 214
rect 3148 206 3154 214
rect 3154 206 3156 214
rect 6156 196 6164 204
rect 716 156 724 164
rect 812 136 820 144
rect 5900 156 5908 164
rect 6028 156 6036 164
rect 6060 136 6068 144
rect 2028 116 2036 124
rect 5420 116 5428 124
rect 5804 116 5812 124
rect 716 96 724 104
rect 1932 96 1940 104
rect 5452 96 5460 104
rect 5644 96 5652 104
rect 5868 96 5876 104
rect 5996 116 6004 124
rect 2700 56 2708 64
rect 3564 56 3572 64
rect 3852 36 3860 44
rect 4172 36 4180 44
rect 2156 16 2164 24
rect 2316 16 2324 24
rect 2604 16 2612 24
rect 4812 16 4820 24
rect 5964 16 5972 24
rect 6156 16 6164 24
rect 1564 6 1566 14
rect 1566 6 1572 14
rect 1580 6 1588 14
rect 1596 6 1602 14
rect 1602 6 1604 14
rect 4636 6 4638 14
rect 4638 6 4644 14
rect 4652 6 4660 14
rect 4668 6 4674 14
rect 4674 6 4676 14
<< metal4 >>
rect 1066 5804 1078 5806
rect 1066 5796 1068 5804
rect 1076 5796 1078 5804
rect 586 5744 598 5746
rect 586 5736 588 5744
rect 596 5736 598 5744
rect 202 5724 214 5726
rect 202 5716 204 5724
rect 212 5716 214 5724
rect 10 5484 22 5486
rect 10 5476 12 5484
rect 20 5476 22 5484
rect 10 5344 22 5476
rect 202 5464 214 5716
rect 202 5456 204 5464
rect 212 5456 214 5464
rect 202 5454 214 5456
rect 458 5544 470 5546
rect 458 5536 460 5544
rect 468 5536 470 5544
rect 10 5336 12 5344
rect 20 5336 22 5344
rect 10 5334 22 5336
rect 394 5444 406 5446
rect 394 5436 396 5444
rect 404 5436 406 5444
rect 394 5304 406 5436
rect 458 5384 470 5536
rect 586 5444 598 5736
rect 1066 5744 1078 5796
rect 1066 5736 1068 5744
rect 1076 5736 1078 5744
rect 906 5724 918 5726
rect 906 5716 908 5724
rect 916 5716 918 5724
rect 586 5436 588 5444
rect 596 5436 598 5444
rect 586 5434 598 5436
rect 618 5464 630 5466
rect 618 5456 620 5464
rect 628 5456 630 5464
rect 458 5376 460 5384
rect 468 5376 470 5384
rect 458 5374 470 5376
rect 394 5296 396 5304
rect 404 5296 406 5304
rect 394 5294 406 5296
rect 618 5284 630 5456
rect 618 5276 620 5284
rect 628 5276 630 5284
rect 618 5274 630 5276
rect 906 5344 918 5716
rect 1034 5444 1046 5446
rect 1034 5436 1036 5444
rect 1044 5436 1046 5444
rect 906 5336 908 5344
rect 916 5336 918 5344
rect 138 5184 150 5186
rect 138 5176 140 5184
rect 148 5176 150 5184
rect 74 5064 86 5066
rect 74 5056 76 5064
rect 84 5056 86 5064
rect 10 4584 22 4586
rect 10 4576 12 4584
rect 20 4576 22 4584
rect 10 4544 22 4576
rect 10 4536 12 4544
rect 20 4536 22 4544
rect 10 4534 22 4536
rect 74 4524 86 5056
rect 74 4516 76 4524
rect 84 4516 86 4524
rect 74 4514 86 4516
rect 106 4664 118 4666
rect 106 4656 108 4664
rect 116 4656 118 4664
rect 42 4484 54 4486
rect 42 4476 44 4484
rect 52 4476 54 4484
rect 42 4344 54 4476
rect 42 4336 44 4344
rect 52 4336 54 4344
rect 10 3964 22 3966
rect 10 3956 12 3964
rect 20 3956 22 3964
rect 10 3884 22 3956
rect 10 3876 12 3884
rect 20 3876 22 3884
rect 10 3874 22 3876
rect 42 3684 54 4336
rect 106 3724 118 4656
rect 138 4644 150 5176
rect 906 5084 918 5336
rect 906 5076 908 5084
rect 916 5076 918 5084
rect 842 4944 854 4946
rect 842 4936 844 4944
rect 852 4936 854 4944
rect 554 4844 566 4846
rect 554 4836 556 4844
rect 564 4836 566 4844
rect 138 4636 140 4644
rect 148 4636 150 4644
rect 138 4634 150 4636
rect 202 4644 214 4646
rect 202 4636 204 4644
rect 212 4636 214 4644
rect 202 4344 214 4636
rect 202 4336 204 4344
rect 212 4336 214 4344
rect 202 4334 214 4336
rect 490 4524 502 4526
rect 490 4516 492 4524
rect 500 4516 502 4524
rect 458 4304 470 4306
rect 458 4296 460 4304
rect 468 4296 470 4304
rect 170 4284 182 4286
rect 170 4276 172 4284
rect 180 4276 182 4284
rect 170 4004 182 4276
rect 170 3996 172 4004
rect 180 3996 182 4004
rect 170 3994 182 3996
rect 330 4284 342 4286
rect 330 4276 332 4284
rect 340 4276 342 4284
rect 330 3824 342 4276
rect 330 3816 332 3824
rect 340 3816 342 3824
rect 330 3814 342 3816
rect 362 4244 374 4246
rect 362 4236 364 4244
rect 372 4236 374 4244
rect 362 4104 374 4236
rect 362 4096 364 4104
rect 372 4096 374 4104
rect 106 3716 108 3724
rect 116 3716 118 3724
rect 106 3714 118 3716
rect 170 3744 182 3746
rect 170 3736 172 3744
rect 180 3736 182 3744
rect 42 3676 44 3684
rect 52 3676 54 3684
rect 42 3674 54 3676
rect 138 3504 150 3506
rect 138 3496 140 3504
rect 148 3496 150 3504
rect 138 3064 150 3496
rect 138 3056 140 3064
rect 148 3056 150 3064
rect 138 3054 150 3056
rect 170 3044 182 3736
rect 266 3684 278 3686
rect 266 3676 268 3684
rect 276 3676 278 3684
rect 234 3404 246 3406
rect 234 3396 236 3404
rect 244 3396 246 3404
rect 234 3344 246 3396
rect 234 3336 236 3344
rect 244 3336 246 3344
rect 234 3334 246 3336
rect 170 3036 172 3044
rect 180 3036 182 3044
rect 170 3034 182 3036
rect 202 3284 214 3286
rect 202 3276 204 3284
rect 212 3276 214 3284
rect 106 2984 118 2986
rect 106 2976 108 2984
rect 116 2976 118 2984
rect 106 2924 118 2976
rect 106 2916 108 2924
rect 116 2916 118 2924
rect 74 2824 86 2826
rect 74 2816 76 2824
rect 84 2816 86 2824
rect 10 2404 22 2406
rect 10 2396 12 2404
rect 20 2396 22 2404
rect 10 1884 22 2396
rect 74 2384 86 2816
rect 106 2444 118 2916
rect 138 2724 150 2726
rect 138 2716 140 2724
rect 148 2716 150 2724
rect 138 2524 150 2716
rect 202 2684 214 3276
rect 266 3164 278 3676
rect 362 3684 374 4096
rect 362 3676 364 3684
rect 372 3676 374 3684
rect 362 3384 374 3676
rect 458 3564 470 4296
rect 490 4104 502 4516
rect 554 4244 566 4836
rect 810 4764 822 4766
rect 810 4756 812 4764
rect 820 4756 822 4764
rect 650 4684 662 4686
rect 650 4676 652 4684
rect 660 4676 662 4684
rect 650 4504 662 4676
rect 650 4496 652 4504
rect 660 4496 662 4504
rect 554 4236 556 4244
rect 564 4236 566 4244
rect 554 4234 566 4236
rect 586 4284 598 4286
rect 586 4276 588 4284
rect 596 4276 598 4284
rect 490 4096 492 4104
rect 500 4096 502 4104
rect 490 4094 502 4096
rect 522 4144 534 4146
rect 522 4136 524 4144
rect 532 4136 534 4144
rect 458 3556 460 3564
rect 468 3556 470 3564
rect 458 3554 470 3556
rect 490 3704 502 3706
rect 490 3696 492 3704
rect 500 3696 502 3704
rect 490 3604 502 3696
rect 490 3596 492 3604
rect 500 3596 502 3604
rect 362 3376 364 3384
rect 372 3376 374 3384
rect 362 3374 374 3376
rect 266 3156 268 3164
rect 276 3156 278 3164
rect 266 3154 278 3156
rect 298 3304 310 3306
rect 298 3296 300 3304
rect 308 3296 310 3304
rect 234 3084 246 3086
rect 234 3076 236 3084
rect 244 3076 246 3084
rect 234 2844 246 3076
rect 234 2836 236 2844
rect 244 2836 246 2844
rect 234 2834 246 2836
rect 298 3024 310 3296
rect 298 3016 300 3024
rect 308 3016 310 3024
rect 202 2676 204 2684
rect 212 2676 214 2684
rect 202 2674 214 2676
rect 138 2516 140 2524
rect 148 2516 150 2524
rect 138 2514 150 2516
rect 106 2436 108 2444
rect 116 2436 118 2444
rect 106 2434 118 2436
rect 74 2376 76 2384
rect 84 2376 86 2384
rect 74 2374 86 2376
rect 106 2384 118 2386
rect 106 2376 108 2384
rect 116 2376 118 2384
rect 106 2104 118 2376
rect 234 2364 246 2366
rect 234 2356 236 2364
rect 244 2356 246 2364
rect 106 2096 108 2104
rect 116 2096 118 2104
rect 106 2094 118 2096
rect 138 2284 150 2286
rect 138 2276 140 2284
rect 148 2276 150 2284
rect 138 2064 150 2276
rect 138 2056 140 2064
rect 148 2056 150 2064
rect 138 2054 150 2056
rect 234 2044 246 2356
rect 234 2036 236 2044
rect 244 2036 246 2044
rect 10 1876 12 1884
rect 20 1876 22 1884
rect 10 1874 22 1876
rect 74 2024 86 2026
rect 74 2016 76 2024
rect 84 2016 86 2024
rect 42 1664 54 1666
rect 42 1656 44 1664
rect 52 1656 54 1664
rect 42 1364 54 1656
rect 42 1356 44 1364
rect 52 1356 54 1364
rect 42 1354 54 1356
rect 74 1064 86 2016
rect 234 1824 246 2036
rect 234 1816 236 1824
rect 244 1816 246 1824
rect 234 1814 246 1816
rect 266 2264 278 2266
rect 266 2256 268 2264
rect 276 2256 278 2264
rect 266 1824 278 2256
rect 298 2264 310 3016
rect 330 3164 342 3166
rect 330 3156 332 3164
rect 340 3156 342 3164
rect 330 3004 342 3156
rect 330 2996 332 3004
rect 340 2996 342 3004
rect 330 2994 342 2996
rect 490 2964 502 3596
rect 522 3244 534 4136
rect 586 4064 598 4276
rect 586 4056 588 4064
rect 596 4056 598 4064
rect 586 4054 598 4056
rect 650 3884 662 4496
rect 682 4484 694 4486
rect 682 4476 684 4484
rect 692 4476 694 4484
rect 682 4264 694 4476
rect 682 4256 684 4264
rect 692 4256 694 4264
rect 682 4254 694 4256
rect 650 3876 652 3884
rect 660 3876 662 3884
rect 650 3874 662 3876
rect 682 3864 694 3866
rect 682 3856 684 3864
rect 692 3856 694 3864
rect 618 3824 630 3826
rect 618 3816 620 3824
rect 628 3816 630 3824
rect 522 3236 524 3244
rect 532 3236 534 3244
rect 522 3234 534 3236
rect 554 3644 566 3646
rect 554 3636 556 3644
rect 564 3636 566 3644
rect 490 2956 492 2964
rect 500 2956 502 2964
rect 490 2954 502 2956
rect 522 3084 534 3086
rect 522 3076 524 3084
rect 532 3076 534 3084
rect 522 2944 534 3076
rect 554 3064 566 3636
rect 554 3056 556 3064
rect 564 3056 566 3064
rect 554 3054 566 3056
rect 586 3344 598 3346
rect 586 3336 588 3344
rect 596 3336 598 3344
rect 522 2936 524 2944
rect 532 2936 534 2944
rect 522 2934 534 2936
rect 554 2904 566 2906
rect 554 2896 556 2904
rect 564 2896 566 2904
rect 362 2824 374 2826
rect 362 2816 364 2824
rect 372 2816 374 2824
rect 362 2484 374 2816
rect 458 2824 470 2826
rect 458 2816 460 2824
rect 468 2816 470 2824
rect 426 2764 438 2766
rect 426 2756 428 2764
rect 436 2756 438 2764
rect 426 2644 438 2756
rect 426 2636 428 2644
rect 436 2636 438 2644
rect 426 2634 438 2636
rect 362 2476 364 2484
rect 372 2476 374 2484
rect 362 2474 374 2476
rect 458 2484 470 2816
rect 522 2584 534 2586
rect 522 2576 524 2584
rect 532 2576 534 2584
rect 522 2544 534 2576
rect 522 2536 524 2544
rect 532 2536 534 2544
rect 522 2534 534 2536
rect 458 2476 460 2484
rect 468 2476 470 2484
rect 458 2474 470 2476
rect 490 2484 502 2486
rect 490 2476 492 2484
rect 500 2476 502 2484
rect 426 2424 438 2426
rect 426 2416 428 2424
rect 436 2416 438 2424
rect 394 2404 406 2406
rect 394 2396 396 2404
rect 404 2396 406 2404
rect 298 2256 300 2264
rect 308 2256 310 2264
rect 298 2004 310 2256
rect 362 2364 374 2366
rect 362 2356 364 2364
rect 372 2356 374 2364
rect 298 1996 300 2004
rect 308 1996 310 2004
rect 298 1994 310 1996
rect 330 2244 342 2246
rect 330 2236 332 2244
rect 340 2236 342 2244
rect 266 1816 268 1824
rect 276 1816 278 1824
rect 266 1814 278 1816
rect 138 1784 150 1786
rect 138 1776 140 1784
rect 148 1776 150 1784
rect 106 1364 118 1366
rect 106 1356 108 1364
rect 116 1356 118 1364
rect 106 1084 118 1356
rect 138 1104 150 1776
rect 330 1724 342 2236
rect 362 1944 374 2356
rect 394 2084 406 2396
rect 426 2304 438 2416
rect 426 2296 428 2304
rect 436 2296 438 2304
rect 426 2294 438 2296
rect 490 2244 502 2476
rect 554 2324 566 2896
rect 586 2764 598 3336
rect 618 3284 630 3816
rect 618 3276 620 3284
rect 628 3276 630 3284
rect 618 3274 630 3276
rect 618 3064 630 3066
rect 618 3056 620 3064
rect 628 3056 630 3064
rect 618 2884 630 3056
rect 618 2876 620 2884
rect 628 2876 630 2884
rect 618 2874 630 2876
rect 650 2924 662 2926
rect 650 2916 652 2924
rect 660 2916 662 2924
rect 586 2756 588 2764
rect 596 2756 598 2764
rect 586 2754 598 2756
rect 650 2724 662 2916
rect 650 2716 652 2724
rect 660 2716 662 2724
rect 650 2714 662 2716
rect 682 2504 694 3856
rect 778 3704 790 3706
rect 778 3696 780 3704
rect 788 3696 790 3704
rect 682 2496 684 2504
rect 692 2496 694 2504
rect 618 2344 630 2346
rect 618 2336 620 2344
rect 628 2336 630 2344
rect 554 2316 556 2324
rect 564 2316 566 2324
rect 554 2314 566 2316
rect 586 2324 598 2326
rect 586 2316 588 2324
rect 596 2316 598 2324
rect 490 2236 492 2244
rect 500 2236 502 2244
rect 490 2234 502 2236
rect 394 2076 396 2084
rect 404 2076 406 2084
rect 394 2074 406 2076
rect 490 2204 502 2206
rect 490 2196 492 2204
rect 500 2196 502 2204
rect 362 1936 364 1944
rect 372 1936 374 1944
rect 362 1934 374 1936
rect 490 1944 502 2196
rect 586 2004 598 2316
rect 586 1996 588 2004
rect 596 1996 598 2004
rect 586 1994 598 1996
rect 618 2004 630 2336
rect 618 1996 620 2004
rect 628 1996 630 2004
rect 618 1994 630 1996
rect 490 1936 492 1944
rect 500 1936 502 1944
rect 490 1934 502 1936
rect 554 1984 566 1986
rect 554 1976 556 1984
rect 564 1976 566 1984
rect 522 1904 534 1906
rect 522 1896 524 1904
rect 532 1896 534 1904
rect 490 1864 502 1866
rect 490 1856 492 1864
rect 500 1856 502 1864
rect 330 1716 332 1724
rect 340 1716 342 1724
rect 330 1714 342 1716
rect 458 1784 470 1786
rect 458 1776 460 1784
rect 468 1776 470 1784
rect 458 1704 470 1776
rect 458 1696 460 1704
rect 468 1696 470 1704
rect 458 1694 470 1696
rect 330 1624 342 1626
rect 330 1616 332 1624
rect 340 1616 342 1624
rect 138 1096 140 1104
rect 148 1096 150 1104
rect 138 1094 150 1096
rect 234 1364 246 1366
rect 234 1356 236 1364
rect 244 1356 246 1364
rect 106 1076 108 1084
rect 116 1076 118 1084
rect 106 1074 118 1076
rect 74 1056 76 1064
rect 84 1056 86 1064
rect 74 1054 86 1056
rect 234 704 246 1356
rect 234 696 236 704
rect 244 696 246 704
rect 234 694 246 696
rect 266 964 278 966
rect 266 956 268 964
rect 276 956 278 964
rect 266 664 278 956
rect 330 964 342 1616
rect 490 1624 502 1856
rect 522 1704 534 1896
rect 522 1696 524 1704
rect 532 1696 534 1704
rect 522 1694 534 1696
rect 490 1616 492 1624
rect 500 1616 502 1624
rect 490 1614 502 1616
rect 522 1624 534 1626
rect 522 1616 524 1624
rect 532 1616 534 1624
rect 522 1504 534 1616
rect 522 1496 524 1504
rect 532 1496 534 1504
rect 522 1494 534 1496
rect 554 1384 566 1976
rect 682 1884 694 2496
rect 682 1876 684 1884
rect 692 1876 694 1884
rect 682 1874 694 1876
rect 714 3644 726 3646
rect 714 3636 716 3644
rect 724 3636 726 3644
rect 714 3444 726 3636
rect 714 3436 716 3444
rect 724 3436 726 3444
rect 714 3344 726 3436
rect 714 3336 716 3344
rect 724 3336 726 3344
rect 714 2684 726 3336
rect 746 3404 758 3406
rect 746 3396 748 3404
rect 756 3396 758 3404
rect 746 3224 758 3396
rect 746 3216 748 3224
rect 756 3216 758 3224
rect 746 3214 758 3216
rect 778 3164 790 3696
rect 778 3156 780 3164
rect 788 3156 790 3164
rect 778 3154 790 3156
rect 714 2676 716 2684
rect 724 2676 726 2684
rect 714 1884 726 2676
rect 714 1876 716 1884
rect 724 1876 726 1884
rect 650 1804 662 1806
rect 650 1796 652 1804
rect 660 1796 662 1804
rect 650 1724 662 1796
rect 650 1716 652 1724
rect 660 1716 662 1724
rect 650 1714 662 1716
rect 682 1724 694 1726
rect 682 1716 684 1724
rect 692 1716 694 1724
rect 650 1624 662 1626
rect 650 1616 652 1624
rect 660 1616 662 1624
rect 554 1376 556 1384
rect 564 1376 566 1384
rect 554 1374 566 1376
rect 586 1424 598 1426
rect 586 1416 588 1424
rect 596 1416 598 1424
rect 586 1324 598 1416
rect 586 1316 588 1324
rect 596 1316 598 1324
rect 586 1314 598 1316
rect 618 1384 630 1386
rect 618 1376 620 1384
rect 628 1376 630 1384
rect 522 1224 534 1226
rect 522 1216 524 1224
rect 532 1216 534 1224
rect 330 956 332 964
rect 340 956 342 964
rect 330 904 342 956
rect 330 896 332 904
rect 340 896 342 904
rect 330 894 342 896
rect 426 1004 438 1006
rect 426 996 428 1004
rect 436 996 438 1004
rect 266 656 268 664
rect 276 656 278 664
rect 266 564 278 656
rect 266 556 268 564
rect 276 556 278 564
rect 266 554 278 556
rect 426 544 438 996
rect 426 536 428 544
rect 436 536 438 544
rect 426 534 438 536
rect 458 624 470 626
rect 458 616 460 624
rect 468 616 470 624
rect 458 364 470 616
rect 522 404 534 1216
rect 618 1164 630 1376
rect 618 1156 620 1164
rect 628 1156 630 1164
rect 618 1154 630 1156
rect 522 396 524 404
rect 532 396 534 404
rect 522 394 534 396
rect 554 504 566 506
rect 554 496 556 504
rect 564 496 566 504
rect 458 356 460 364
rect 468 356 470 364
rect 458 354 470 356
rect 554 284 566 496
rect 650 504 662 1616
rect 682 1604 694 1716
rect 682 1596 684 1604
rect 692 1596 694 1604
rect 682 1594 694 1596
rect 714 1524 726 1876
rect 714 1516 716 1524
rect 724 1516 726 1524
rect 714 1124 726 1516
rect 746 2964 758 2966
rect 746 2956 748 2964
rect 756 2956 758 2964
rect 746 2304 758 2956
rect 778 2744 790 2746
rect 778 2736 780 2744
rect 788 2736 790 2744
rect 778 2544 790 2736
rect 810 2724 822 4756
rect 842 4144 854 4936
rect 842 4136 844 4144
rect 852 4136 854 4144
rect 842 4134 854 4136
rect 906 4664 918 5076
rect 970 5404 982 5406
rect 970 5396 972 5404
rect 980 5396 982 5404
rect 970 4944 982 5396
rect 970 4936 972 4944
rect 980 4936 982 4944
rect 970 4764 982 4936
rect 1034 4944 1046 5436
rect 1034 4936 1036 4944
rect 1044 4936 1046 4944
rect 1034 4934 1046 4936
rect 1066 5284 1078 5736
rect 1130 5804 1142 5806
rect 1130 5796 1132 5804
rect 1140 5796 1142 5804
rect 1130 5644 1142 5796
rect 1130 5636 1132 5644
rect 1140 5636 1142 5644
rect 1130 5634 1142 5636
rect 1450 5684 1462 5686
rect 1450 5676 1452 5684
rect 1460 5676 1462 5684
rect 1258 5524 1270 5526
rect 1258 5516 1260 5524
rect 1268 5516 1270 5524
rect 1258 5384 1270 5516
rect 1258 5376 1260 5384
rect 1268 5376 1270 5384
rect 1258 5374 1270 5376
rect 1354 5524 1366 5526
rect 1354 5516 1356 5524
rect 1364 5516 1366 5524
rect 1066 5276 1068 5284
rect 1076 5276 1078 5284
rect 970 4756 972 4764
rect 980 4756 982 4764
rect 970 4754 982 4756
rect 906 4656 908 4664
rect 916 4656 918 4664
rect 842 4104 854 4106
rect 842 4096 844 4104
rect 852 4096 854 4104
rect 842 3784 854 4096
rect 842 3776 844 3784
rect 852 3776 854 3784
rect 842 3774 854 3776
rect 810 2716 812 2724
rect 820 2716 822 2724
rect 810 2714 822 2716
rect 842 3724 854 3726
rect 842 3716 844 3724
rect 852 3716 854 3724
rect 778 2536 780 2544
rect 788 2536 790 2544
rect 778 2534 790 2536
rect 842 2544 854 3716
rect 874 3704 886 3706
rect 874 3696 876 3704
rect 884 3696 886 3704
rect 874 3364 886 3696
rect 874 3356 876 3364
rect 884 3356 886 3364
rect 874 3354 886 3356
rect 906 3344 918 4656
rect 938 4644 950 4646
rect 938 4636 940 4644
rect 948 4636 950 4644
rect 938 4104 950 4636
rect 1034 4584 1046 4586
rect 1034 4576 1036 4584
rect 1044 4576 1046 4584
rect 1034 4364 1046 4576
rect 1034 4356 1036 4364
rect 1044 4356 1046 4364
rect 1034 4354 1046 4356
rect 938 4096 940 4104
rect 948 4096 950 4104
rect 938 4094 950 4096
rect 1034 3884 1046 3886
rect 1034 3876 1036 3884
rect 1044 3876 1046 3884
rect 938 3644 950 3646
rect 938 3636 940 3644
rect 948 3636 950 3644
rect 938 3424 950 3636
rect 938 3416 940 3424
rect 948 3416 950 3424
rect 938 3414 950 3416
rect 1034 3364 1046 3876
rect 1034 3356 1036 3364
rect 1044 3356 1046 3364
rect 1034 3354 1046 3356
rect 906 3336 908 3344
rect 916 3336 918 3344
rect 874 3164 886 3166
rect 874 3156 876 3164
rect 884 3156 886 3164
rect 874 3044 886 3156
rect 874 3036 876 3044
rect 884 3036 886 3044
rect 874 3034 886 3036
rect 842 2536 844 2544
rect 852 2536 854 2544
rect 746 2296 748 2304
rect 756 2296 758 2304
rect 746 2104 758 2296
rect 746 2096 748 2104
rect 756 2096 758 2104
rect 746 1324 758 2096
rect 842 1904 854 2536
rect 842 1896 844 1904
rect 852 1896 854 1904
rect 842 1894 854 1896
rect 874 2084 886 2086
rect 874 2076 876 2084
rect 884 2076 886 2084
rect 810 1844 822 1846
rect 810 1836 812 1844
rect 820 1836 822 1844
rect 778 1524 790 1526
rect 778 1516 780 1524
rect 788 1516 790 1524
rect 778 1344 790 1516
rect 810 1524 822 1836
rect 842 1744 854 1746
rect 842 1736 844 1744
rect 852 1736 854 1744
rect 842 1584 854 1736
rect 842 1576 844 1584
rect 852 1576 854 1584
rect 842 1574 854 1576
rect 810 1516 812 1524
rect 820 1516 822 1524
rect 810 1514 822 1516
rect 842 1384 854 1386
rect 842 1376 844 1384
rect 852 1376 854 1384
rect 778 1336 780 1344
rect 788 1336 790 1344
rect 778 1334 790 1336
rect 810 1344 822 1346
rect 810 1336 812 1344
rect 820 1336 822 1344
rect 746 1316 748 1324
rect 756 1316 758 1324
rect 746 1314 758 1316
rect 714 1116 716 1124
rect 724 1116 726 1124
rect 714 1114 726 1116
rect 810 1084 822 1336
rect 842 1304 854 1376
rect 842 1296 844 1304
rect 852 1296 854 1304
rect 842 1294 854 1296
rect 874 1184 886 2076
rect 906 1924 918 3336
rect 1002 3324 1014 3326
rect 1002 3316 1004 3324
rect 1012 3316 1014 3324
rect 938 3284 950 3286
rect 938 3276 940 3284
rect 948 3276 950 3284
rect 938 2944 950 3276
rect 1002 3064 1014 3316
rect 1066 3324 1078 5276
rect 1354 5264 1366 5516
rect 1450 5524 1462 5676
rect 1450 5516 1452 5524
rect 1460 5516 1462 5524
rect 1450 5514 1462 5516
rect 1560 5614 1608 5840
rect 3112 5814 3160 5840
rect 3112 5806 3116 5814
rect 3124 5806 3132 5814
rect 3140 5806 3148 5814
rect 3156 5806 3160 5814
rect 3050 5804 3062 5806
rect 3050 5796 3052 5804
rect 3060 5796 3062 5804
rect 1962 5764 1974 5766
rect 1962 5756 1964 5764
rect 1972 5756 1974 5764
rect 1962 5726 1974 5756
rect 1962 5724 2038 5726
rect 1962 5716 2028 5724
rect 2036 5716 2038 5724
rect 1962 5714 2038 5716
rect 1560 5606 1564 5614
rect 1572 5606 1580 5614
rect 1588 5606 1596 5614
rect 1604 5606 1608 5614
rect 1514 5464 1526 5466
rect 1514 5456 1516 5464
rect 1524 5456 1526 5464
rect 1354 5256 1356 5264
rect 1364 5256 1366 5264
rect 1354 5254 1366 5256
rect 1418 5424 1430 5426
rect 1418 5416 1420 5424
rect 1428 5416 1430 5424
rect 1418 5344 1430 5416
rect 1418 5336 1420 5344
rect 1428 5336 1430 5344
rect 1418 5084 1430 5336
rect 1418 5076 1420 5084
rect 1428 5076 1430 5084
rect 1258 5004 1270 5006
rect 1258 4996 1260 5004
rect 1268 4996 1270 5004
rect 1194 4804 1206 4806
rect 1194 4796 1196 4804
rect 1204 4796 1206 4804
rect 1098 4264 1110 4266
rect 1098 4256 1100 4264
rect 1108 4256 1110 4264
rect 1098 3864 1110 4256
rect 1194 4244 1206 4796
rect 1194 4236 1196 4244
rect 1204 4236 1206 4244
rect 1194 4234 1206 4236
rect 1130 4204 1142 4206
rect 1130 4196 1132 4204
rect 1140 4196 1142 4204
rect 1130 4124 1142 4196
rect 1130 4116 1132 4124
rect 1140 4116 1142 4124
rect 1130 4114 1142 4116
rect 1098 3856 1100 3864
rect 1108 3856 1110 3864
rect 1098 3854 1110 3856
rect 1162 3884 1174 3886
rect 1162 3876 1164 3884
rect 1172 3876 1174 3884
rect 1130 3844 1142 3846
rect 1130 3836 1132 3844
rect 1140 3836 1142 3844
rect 1130 3704 1142 3836
rect 1130 3696 1132 3704
rect 1140 3696 1142 3704
rect 1066 3316 1068 3324
rect 1076 3316 1078 3324
rect 1066 3314 1078 3316
rect 1098 3324 1110 3326
rect 1098 3316 1100 3324
rect 1108 3316 1110 3324
rect 1002 3056 1004 3064
rect 1012 3056 1014 3064
rect 1002 3054 1014 3056
rect 1066 3204 1078 3206
rect 1066 3196 1068 3204
rect 1076 3196 1078 3204
rect 1066 3064 1078 3196
rect 1066 3056 1068 3064
rect 1076 3056 1078 3064
rect 1066 3054 1078 3056
rect 938 2936 940 2944
rect 948 2936 950 2944
rect 938 2934 950 2936
rect 1066 2944 1078 2946
rect 1066 2936 1068 2944
rect 1076 2936 1078 2944
rect 938 2884 950 2886
rect 938 2876 940 2884
rect 948 2876 950 2884
rect 938 2604 950 2876
rect 1034 2864 1046 2866
rect 1034 2856 1036 2864
rect 1044 2856 1046 2864
rect 938 2596 940 2604
rect 948 2596 950 2604
rect 938 2594 950 2596
rect 970 2744 982 2746
rect 970 2736 972 2744
rect 980 2736 982 2744
rect 906 1916 908 1924
rect 916 1916 918 1924
rect 906 1914 918 1916
rect 970 2484 982 2736
rect 970 2476 972 2484
rect 980 2476 982 2484
rect 906 1824 918 1826
rect 906 1816 908 1824
rect 916 1816 918 1824
rect 906 1744 918 1816
rect 906 1736 908 1744
rect 916 1736 918 1744
rect 906 1734 918 1736
rect 938 1804 950 1806
rect 938 1796 940 1804
rect 948 1796 950 1804
rect 938 1484 950 1796
rect 938 1476 940 1484
rect 948 1476 950 1484
rect 938 1474 950 1476
rect 970 1624 982 2476
rect 1002 2624 1014 2626
rect 1002 2616 1004 2624
rect 1012 2616 1014 2624
rect 1002 2244 1014 2616
rect 1002 2236 1004 2244
rect 1012 2236 1014 2244
rect 1002 2234 1014 2236
rect 970 1616 972 1624
rect 980 1616 982 1624
rect 970 1464 982 1616
rect 970 1456 972 1464
rect 980 1456 982 1464
rect 970 1454 982 1456
rect 1034 1824 1046 2856
rect 1066 2564 1078 2936
rect 1066 2556 1068 2564
rect 1076 2556 1078 2564
rect 1066 2554 1078 2556
rect 1098 2684 1110 3316
rect 1130 3204 1142 3696
rect 1162 3664 1174 3876
rect 1162 3656 1164 3664
rect 1172 3656 1174 3664
rect 1162 3654 1174 3656
rect 1226 3664 1238 3666
rect 1226 3656 1228 3664
rect 1236 3656 1238 3664
rect 1130 3196 1132 3204
rect 1140 3196 1142 3204
rect 1130 3194 1142 3196
rect 1194 3444 1206 3446
rect 1194 3436 1196 3444
rect 1204 3436 1206 3444
rect 1162 3004 1174 3006
rect 1162 2996 1164 3004
rect 1172 2996 1174 3004
rect 1162 2924 1174 2996
rect 1162 2916 1164 2924
rect 1172 2916 1174 2924
rect 1162 2914 1174 2916
rect 1098 2676 1100 2684
rect 1108 2676 1110 2684
rect 1034 1816 1036 1824
rect 1044 1816 1046 1824
rect 1034 1524 1046 1816
rect 1034 1516 1036 1524
rect 1044 1516 1046 1524
rect 1002 1404 1014 1406
rect 1002 1396 1004 1404
rect 1012 1396 1014 1404
rect 970 1384 982 1386
rect 970 1376 972 1384
rect 980 1376 982 1384
rect 970 1324 982 1376
rect 970 1316 972 1324
rect 980 1316 982 1324
rect 970 1314 982 1316
rect 1002 1304 1014 1396
rect 1034 1344 1046 1516
rect 1066 2424 1078 2426
rect 1066 2416 1068 2424
rect 1076 2416 1078 2424
rect 1066 1744 1078 2416
rect 1066 1736 1068 1744
rect 1076 1736 1078 1744
rect 1066 1484 1078 1736
rect 1098 1684 1110 2676
rect 1162 2844 1174 2846
rect 1162 2836 1164 2844
rect 1172 2836 1174 2844
rect 1130 2664 1142 2666
rect 1130 2656 1132 2664
rect 1140 2656 1142 2664
rect 1130 2324 1142 2656
rect 1162 2604 1174 2836
rect 1162 2596 1164 2604
rect 1172 2596 1174 2604
rect 1162 2594 1174 2596
rect 1130 2316 1132 2324
rect 1140 2316 1142 2324
rect 1130 2314 1142 2316
rect 1194 2584 1206 3436
rect 1226 3304 1238 3656
rect 1226 3296 1228 3304
rect 1236 3296 1238 3304
rect 1226 2724 1238 3296
rect 1226 2716 1228 2724
rect 1236 2716 1238 2724
rect 1226 2714 1238 2716
rect 1258 3624 1270 4996
rect 1386 4764 1398 4766
rect 1386 4756 1388 4764
rect 1396 4756 1398 4764
rect 1290 4644 1302 4646
rect 1290 4636 1292 4644
rect 1300 4636 1302 4644
rect 1290 4164 1302 4636
rect 1290 4156 1292 4164
rect 1300 4156 1302 4164
rect 1290 4154 1302 4156
rect 1354 4164 1366 4166
rect 1354 4156 1356 4164
rect 1364 4156 1366 4164
rect 1322 3884 1334 3886
rect 1322 3876 1324 3884
rect 1332 3876 1334 3884
rect 1322 3824 1334 3876
rect 1322 3816 1324 3824
rect 1332 3816 1334 3824
rect 1258 3616 1260 3624
rect 1268 3616 1270 3624
rect 1194 2576 1196 2584
rect 1204 2576 1206 2584
rect 1130 2284 1142 2286
rect 1130 2276 1132 2284
rect 1140 2276 1142 2284
rect 1130 2044 1142 2276
rect 1130 2036 1132 2044
rect 1140 2036 1142 2044
rect 1130 2034 1142 2036
rect 1162 1964 1174 1966
rect 1162 1956 1164 1964
rect 1172 1956 1174 1964
rect 1162 1924 1174 1956
rect 1162 1916 1164 1924
rect 1172 1916 1174 1924
rect 1162 1914 1174 1916
rect 1162 1784 1174 1786
rect 1162 1776 1164 1784
rect 1172 1776 1174 1784
rect 1098 1676 1100 1684
rect 1108 1676 1110 1684
rect 1098 1674 1110 1676
rect 1130 1724 1142 1726
rect 1130 1716 1132 1724
rect 1140 1716 1142 1724
rect 1066 1476 1068 1484
rect 1076 1476 1078 1484
rect 1066 1474 1078 1476
rect 1034 1336 1036 1344
rect 1044 1336 1046 1344
rect 1034 1334 1046 1336
rect 1002 1296 1004 1304
rect 1012 1296 1014 1304
rect 1002 1294 1014 1296
rect 1130 1204 1142 1716
rect 1162 1664 1174 1776
rect 1162 1656 1164 1664
rect 1172 1656 1174 1664
rect 1162 1654 1174 1656
rect 1194 1504 1206 2576
rect 1258 2704 1270 3616
rect 1290 3744 1302 3746
rect 1290 3736 1292 3744
rect 1300 3736 1302 3744
rect 1290 3344 1302 3736
rect 1290 3336 1292 3344
rect 1300 3336 1302 3344
rect 1290 3334 1302 3336
rect 1322 3704 1334 3816
rect 1354 3724 1366 4156
rect 1386 4104 1398 4756
rect 1386 4096 1388 4104
rect 1396 4096 1398 4104
rect 1386 4094 1398 4096
rect 1354 3716 1356 3724
rect 1364 3716 1366 3724
rect 1354 3714 1366 3716
rect 1418 3784 1430 5076
rect 1418 3776 1420 3784
rect 1428 3776 1430 3784
rect 1322 3696 1324 3704
rect 1332 3696 1334 3704
rect 1258 2696 1260 2704
rect 1268 2696 1270 2704
rect 1226 2564 1238 2566
rect 1226 2556 1228 2564
rect 1236 2556 1238 2564
rect 1226 2504 1238 2556
rect 1226 2496 1228 2504
rect 1236 2496 1238 2504
rect 1226 2494 1238 2496
rect 1258 1764 1270 2696
rect 1258 1756 1260 1764
rect 1268 1756 1270 1764
rect 1258 1754 1270 1756
rect 1290 3224 1302 3226
rect 1290 3216 1292 3224
rect 1300 3216 1302 3224
rect 1290 1724 1302 3216
rect 1322 2964 1334 3696
rect 1354 3684 1366 3686
rect 1354 3676 1356 3684
rect 1364 3676 1366 3684
rect 1354 3564 1366 3676
rect 1354 3556 1356 3564
rect 1364 3556 1366 3564
rect 1354 3554 1366 3556
rect 1386 3684 1398 3686
rect 1386 3676 1388 3684
rect 1396 3676 1398 3684
rect 1322 2956 1324 2964
rect 1332 2956 1334 2964
rect 1322 2544 1334 2956
rect 1386 3304 1398 3676
rect 1386 3296 1388 3304
rect 1396 3296 1398 3304
rect 1386 2744 1398 3296
rect 1386 2736 1388 2744
rect 1396 2736 1398 2744
rect 1386 2734 1398 2736
rect 1418 2844 1430 3776
rect 1450 3724 1462 3726
rect 1450 3716 1452 3724
rect 1460 3716 1462 3724
rect 1450 3324 1462 3716
rect 1450 3316 1452 3324
rect 1460 3316 1462 3324
rect 1450 3314 1462 3316
rect 1482 3404 1494 3406
rect 1482 3396 1484 3404
rect 1492 3396 1494 3404
rect 1482 3324 1494 3396
rect 1482 3316 1484 3324
rect 1492 3316 1494 3324
rect 1482 3314 1494 3316
rect 1450 3204 1462 3206
rect 1450 3196 1452 3204
rect 1460 3196 1462 3204
rect 1450 3044 1462 3196
rect 1450 3036 1452 3044
rect 1460 3036 1462 3044
rect 1450 3034 1462 3036
rect 1418 2836 1420 2844
rect 1428 2836 1430 2844
rect 1418 2744 1430 2836
rect 1418 2736 1420 2744
rect 1428 2736 1430 2744
rect 1418 2734 1430 2736
rect 1514 2944 1526 5456
rect 1514 2936 1516 2944
rect 1524 2936 1526 2944
rect 1322 2536 1324 2544
rect 1332 2536 1334 2544
rect 1322 2534 1334 2536
rect 1354 2604 1366 2606
rect 1354 2596 1356 2604
rect 1364 2596 1366 2604
rect 1354 2324 1366 2596
rect 1514 2524 1526 2936
rect 1514 2516 1516 2524
rect 1524 2516 1526 2524
rect 1418 2464 1430 2466
rect 1418 2456 1420 2464
rect 1428 2456 1430 2464
rect 1354 2316 1356 2324
rect 1364 2316 1366 2324
rect 1354 2314 1366 2316
rect 1386 2384 1398 2386
rect 1386 2376 1388 2384
rect 1396 2376 1398 2384
rect 1386 1784 1398 2376
rect 1418 2284 1430 2456
rect 1418 2276 1420 2284
rect 1428 2276 1430 2284
rect 1418 2274 1430 2276
rect 1514 2304 1526 2516
rect 1514 2296 1516 2304
rect 1524 2296 1526 2304
rect 1482 2004 1494 2006
rect 1482 1996 1484 2004
rect 1492 1996 1494 2004
rect 1482 1844 1494 1996
rect 1482 1836 1484 1844
rect 1492 1836 1494 1844
rect 1482 1834 1494 1836
rect 1386 1776 1388 1784
rect 1396 1776 1398 1784
rect 1386 1774 1398 1776
rect 1290 1716 1292 1724
rect 1300 1716 1302 1724
rect 1290 1714 1302 1716
rect 1514 1644 1526 2296
rect 1514 1636 1516 1644
rect 1524 1636 1526 1644
rect 1514 1634 1526 1636
rect 1560 5214 1608 5606
rect 1560 5206 1564 5214
rect 1572 5206 1580 5214
rect 1588 5206 1596 5214
rect 1604 5206 1608 5214
rect 1560 4814 1608 5206
rect 2250 5704 2262 5706
rect 2250 5696 2252 5704
rect 2260 5696 2262 5704
rect 1560 4806 1564 4814
rect 1572 4806 1580 4814
rect 1588 4806 1596 4814
rect 1604 4806 1608 4814
rect 1560 4414 1608 4806
rect 1560 4406 1564 4414
rect 1572 4406 1580 4414
rect 1588 4406 1596 4414
rect 1604 4406 1608 4414
rect 1560 4014 1608 4406
rect 1674 5004 1686 5006
rect 1674 4996 1676 5004
rect 1684 4996 1686 5004
rect 1560 4006 1564 4014
rect 1572 4006 1580 4014
rect 1588 4006 1596 4014
rect 1604 4006 1608 4014
rect 1560 3614 1608 4006
rect 1642 4364 1654 4366
rect 1642 4356 1644 4364
rect 1652 4356 1654 4364
rect 1642 3664 1654 4356
rect 1642 3656 1644 3664
rect 1652 3656 1654 3664
rect 1642 3654 1654 3656
rect 1560 3606 1564 3614
rect 1572 3606 1580 3614
rect 1588 3606 1596 3614
rect 1604 3606 1608 3614
rect 1560 3214 1608 3606
rect 1560 3206 1564 3214
rect 1572 3206 1580 3214
rect 1588 3206 1596 3214
rect 1604 3206 1608 3214
rect 1560 2814 1608 3206
rect 1560 2806 1564 2814
rect 1572 2806 1580 2814
rect 1588 2806 1596 2814
rect 1604 2806 1608 2814
rect 1560 2414 1608 2806
rect 1642 3524 1654 3526
rect 1642 3516 1644 3524
rect 1652 3516 1654 3524
rect 1642 3284 1654 3516
rect 1642 3276 1644 3284
rect 1652 3276 1654 3284
rect 1642 2764 1654 3276
rect 1674 3264 1686 4996
rect 1802 5004 1814 5006
rect 1802 4996 1804 5004
rect 1812 4996 1814 5004
rect 1802 3604 1814 4996
rect 2026 4684 2038 4686
rect 2026 4676 2028 4684
rect 2036 4676 2038 4684
rect 2026 3984 2038 4676
rect 2218 4304 2230 4306
rect 2218 4296 2220 4304
rect 2228 4296 2230 4304
rect 2218 4264 2230 4296
rect 2218 4256 2220 4264
rect 2228 4256 2230 4264
rect 2218 4254 2230 4256
rect 2250 4164 2262 5696
rect 2794 5544 2806 5546
rect 2794 5536 2796 5544
rect 2804 5536 2806 5544
rect 2378 5484 2390 5486
rect 2378 5476 2380 5484
rect 2388 5476 2390 5484
rect 2282 5364 2294 5366
rect 2282 5356 2284 5364
rect 2292 5356 2294 5364
rect 2282 5244 2294 5356
rect 2282 5236 2284 5244
rect 2292 5236 2294 5244
rect 2282 5234 2294 5236
rect 2378 4764 2390 5476
rect 2698 5484 2710 5486
rect 2698 5476 2700 5484
rect 2708 5476 2710 5484
rect 2698 5284 2710 5476
rect 2698 5276 2700 5284
rect 2708 5276 2710 5284
rect 2698 5274 2710 5276
rect 2794 5284 2806 5536
rect 2794 5276 2796 5284
rect 2804 5276 2806 5284
rect 2794 5274 2806 5276
rect 2634 5064 2646 5066
rect 2634 5056 2636 5064
rect 2644 5056 2646 5064
rect 2506 5024 2518 5026
rect 2506 5016 2508 5024
rect 2516 5016 2518 5024
rect 2506 4924 2518 5016
rect 2506 4916 2508 4924
rect 2516 4916 2518 4924
rect 2506 4914 2518 4916
rect 2378 4756 2380 4764
rect 2388 4756 2390 4764
rect 2378 4754 2390 4756
rect 2634 4664 2646 5056
rect 3050 4904 3062 5796
rect 3112 5414 3160 5806
rect 4632 5614 4680 5840
rect 5898 5744 5910 5746
rect 5898 5736 5900 5744
rect 5908 5736 5910 5744
rect 4632 5606 4636 5614
rect 4644 5606 4652 5614
rect 4660 5606 4668 5614
rect 4676 5606 4680 5614
rect 3112 5406 3116 5414
rect 3124 5406 3132 5414
rect 3140 5406 3148 5414
rect 3156 5406 3160 5414
rect 3112 5014 3160 5406
rect 3722 5604 3734 5606
rect 3722 5596 3724 5604
rect 3732 5596 3734 5604
rect 3562 5384 3574 5386
rect 3562 5376 3564 5384
rect 3572 5376 3574 5384
rect 3498 5344 3510 5346
rect 3498 5336 3500 5344
rect 3508 5336 3510 5344
rect 3112 5006 3116 5014
rect 3124 5006 3132 5014
rect 3140 5006 3148 5014
rect 3156 5006 3160 5014
rect 3050 4896 3052 4904
rect 3060 4896 3062 4904
rect 3050 4894 3062 4896
rect 3082 4944 3094 4946
rect 3082 4936 3084 4944
rect 3092 4936 3094 4944
rect 3050 4764 3062 4766
rect 3050 4756 3052 4764
rect 3060 4756 3062 4764
rect 2634 4656 2636 4664
rect 2644 4656 2646 4664
rect 2634 4654 2646 4656
rect 2730 4724 2742 4726
rect 2730 4716 2732 4724
rect 2740 4716 2742 4724
rect 2474 4484 2486 4486
rect 2474 4476 2476 4484
rect 2484 4476 2486 4484
rect 2250 4156 2252 4164
rect 2260 4156 2262 4164
rect 2250 4154 2262 4156
rect 2378 4464 2390 4466
rect 2378 4456 2380 4464
rect 2388 4456 2390 4464
rect 2378 4164 2390 4456
rect 2378 4156 2380 4164
rect 2388 4156 2390 4164
rect 2378 4154 2390 4156
rect 2026 3976 2028 3984
rect 2036 3976 2038 3984
rect 2026 3974 2038 3976
rect 2250 4124 2262 4126
rect 2250 4116 2252 4124
rect 2260 4116 2262 4124
rect 1834 3844 1846 3846
rect 1834 3836 1836 3844
rect 1844 3836 1846 3844
rect 1834 3644 1846 3836
rect 2250 3824 2262 4116
rect 2250 3816 2252 3824
rect 2260 3816 2262 3824
rect 2250 3814 2262 3816
rect 1834 3636 1836 3644
rect 1844 3636 1846 3644
rect 1834 3634 1846 3636
rect 2474 3624 2486 4476
rect 2730 4484 2742 4716
rect 2730 4476 2732 4484
rect 2740 4476 2742 4484
rect 2730 4474 2742 4476
rect 3050 4484 3062 4756
rect 3082 4504 3094 4936
rect 3082 4496 3084 4504
rect 3092 4496 3094 4504
rect 3082 4494 3094 4496
rect 3112 4614 3160 5006
rect 3466 5124 3478 5126
rect 3466 5116 3468 5124
rect 3476 5116 3478 5124
rect 3402 4944 3414 4946
rect 3402 4936 3404 4944
rect 3412 4936 3414 4944
rect 3112 4606 3116 4614
rect 3124 4606 3132 4614
rect 3140 4606 3148 4614
rect 3156 4606 3160 4614
rect 3050 4476 3052 4484
rect 3060 4476 3062 4484
rect 3050 4474 3062 4476
rect 2890 4464 2902 4466
rect 2890 4456 2892 4464
rect 2900 4456 2902 4464
rect 2666 4264 2678 4266
rect 2666 4256 2668 4264
rect 2676 4256 2678 4264
rect 2666 4104 2678 4256
rect 2666 4096 2668 4104
rect 2676 4096 2678 4104
rect 2602 4064 2614 4066
rect 2602 4056 2604 4064
rect 2612 4056 2614 4064
rect 2602 3844 2614 4056
rect 2602 3836 2604 3844
rect 2612 3836 2614 3844
rect 2602 3834 2614 3836
rect 2634 3884 2646 3886
rect 2634 3876 2636 3884
rect 2644 3876 2646 3884
rect 2634 3764 2646 3876
rect 2634 3756 2636 3764
rect 2644 3756 2646 3764
rect 2634 3754 2646 3756
rect 2474 3616 2476 3624
rect 2484 3616 2486 3624
rect 2474 3614 2486 3616
rect 2602 3744 2614 3746
rect 2602 3736 2604 3744
rect 2612 3736 2614 3744
rect 1802 3596 1804 3604
rect 1812 3596 1814 3604
rect 1802 3594 1814 3596
rect 2602 3584 2614 3736
rect 2602 3576 2604 3584
rect 2612 3576 2614 3584
rect 2314 3564 2326 3566
rect 2314 3556 2316 3564
rect 2324 3556 2326 3564
rect 2250 3524 2262 3526
rect 2250 3516 2252 3524
rect 2260 3516 2262 3524
rect 1818 3484 1974 3486
rect 1818 3476 1820 3484
rect 1828 3476 1964 3484
rect 1972 3476 1974 3484
rect 1818 3474 1974 3476
rect 2250 3444 2262 3516
rect 2250 3436 2252 3444
rect 2260 3436 2262 3444
rect 2250 3434 2262 3436
rect 2314 3404 2326 3556
rect 2602 3424 2614 3576
rect 2666 3444 2678 4096
rect 2890 4104 2902 4456
rect 2986 4344 2998 4346
rect 2986 4336 2988 4344
rect 2996 4336 2998 4344
rect 2890 4096 2892 4104
rect 2900 4096 2902 4104
rect 2890 4094 2902 4096
rect 2954 4304 2966 4306
rect 2954 4296 2956 4304
rect 2964 4296 2966 4304
rect 2954 4104 2966 4296
rect 2954 4096 2956 4104
rect 2964 4096 2966 4104
rect 2954 4094 2966 4096
rect 2986 4064 2998 4336
rect 2986 4056 2988 4064
rect 2996 4056 2998 4064
rect 2986 4054 2998 4056
rect 3112 4214 3160 4606
rect 3370 4904 3382 4906
rect 3370 4896 3372 4904
rect 3380 4896 3382 4904
rect 3274 4484 3286 4486
rect 3274 4476 3276 4484
rect 3284 4476 3286 4484
rect 3274 4304 3286 4476
rect 3370 4464 3382 4896
rect 3370 4456 3372 4464
rect 3380 4456 3382 4464
rect 3370 4454 3382 4456
rect 3274 4296 3276 4304
rect 3284 4296 3286 4304
rect 3274 4294 3286 4296
rect 3370 4384 3382 4386
rect 3370 4376 3372 4384
rect 3380 4376 3382 4384
rect 3112 4206 3116 4214
rect 3124 4206 3132 4214
rect 3140 4206 3148 4214
rect 3156 4206 3160 4214
rect 3112 3814 3160 4206
rect 3274 4164 3286 4166
rect 3274 4156 3276 4164
rect 3284 4156 3286 4164
rect 3210 3864 3222 3866
rect 3210 3856 3212 3864
rect 3220 3856 3222 3864
rect 3112 3806 3116 3814
rect 3124 3806 3132 3814
rect 3140 3806 3148 3814
rect 3156 3806 3160 3814
rect 3082 3804 3094 3806
rect 3082 3796 3084 3804
rect 3092 3796 3094 3804
rect 3050 3724 3062 3726
rect 3050 3716 3052 3724
rect 3060 3716 3062 3724
rect 2666 3436 2668 3444
rect 2676 3436 2678 3444
rect 2666 3434 2678 3436
rect 2858 3644 2870 3646
rect 2858 3636 2860 3644
rect 2868 3636 2870 3644
rect 2602 3416 2604 3424
rect 2612 3416 2614 3424
rect 2602 3414 2614 3416
rect 2314 3396 2316 3404
rect 2324 3396 2326 3404
rect 2314 3394 2326 3396
rect 1674 3256 1676 3264
rect 1684 3256 1686 3264
rect 1674 3254 1686 3256
rect 1738 3384 1750 3386
rect 1738 3376 1740 3384
rect 1748 3376 1750 3384
rect 1642 2756 1644 2764
rect 1652 2756 1654 2764
rect 1642 2754 1654 2756
rect 1706 2844 1718 2846
rect 1706 2836 1708 2844
rect 1716 2836 1718 2844
rect 1706 2684 1718 2836
rect 1706 2676 1708 2684
rect 1716 2676 1718 2684
rect 1706 2484 1718 2676
rect 1706 2476 1708 2484
rect 1716 2476 1718 2484
rect 1706 2474 1718 2476
rect 1738 2464 1750 3376
rect 1866 3364 1878 3366
rect 1866 3356 1868 3364
rect 1876 3356 1878 3364
rect 1770 3164 1782 3166
rect 1770 3156 1772 3164
rect 1780 3156 1782 3164
rect 1770 2784 1782 3156
rect 1834 3124 1846 3126
rect 1834 3116 1836 3124
rect 1844 3116 1846 3124
rect 1834 2964 1846 3116
rect 1834 2956 1836 2964
rect 1844 2956 1846 2964
rect 1834 2954 1846 2956
rect 1770 2776 1772 2784
rect 1780 2776 1782 2784
rect 1770 2774 1782 2776
rect 1738 2456 1740 2464
rect 1748 2456 1750 2464
rect 1738 2454 1750 2456
rect 1560 2406 1564 2414
rect 1572 2406 1580 2414
rect 1588 2406 1596 2414
rect 1604 2406 1608 2414
rect 1560 2014 1608 2406
rect 1674 2364 1686 2366
rect 1674 2356 1676 2364
rect 1684 2356 1686 2364
rect 1642 2124 1654 2126
rect 1642 2116 1644 2124
rect 1652 2116 1654 2124
rect 1642 2064 1654 2116
rect 1642 2056 1644 2064
rect 1652 2056 1654 2064
rect 1642 2054 1654 2056
rect 1560 2006 1564 2014
rect 1572 2006 1580 2014
rect 1588 2006 1596 2014
rect 1604 2006 1608 2014
rect 1560 1614 1608 2006
rect 1560 1606 1564 1614
rect 1572 1606 1580 1614
rect 1588 1606 1596 1614
rect 1604 1606 1608 1614
rect 1194 1496 1196 1504
rect 1204 1496 1206 1504
rect 1194 1494 1206 1496
rect 1226 1544 1238 1546
rect 1226 1536 1228 1544
rect 1236 1536 1238 1544
rect 1226 1484 1238 1536
rect 1226 1476 1228 1484
rect 1236 1476 1238 1484
rect 1226 1474 1238 1476
rect 1450 1504 1462 1506
rect 1450 1496 1452 1504
rect 1460 1496 1462 1504
rect 1290 1464 1302 1466
rect 1290 1456 1292 1464
rect 1300 1456 1302 1464
rect 1130 1196 1132 1204
rect 1140 1196 1142 1204
rect 1130 1194 1142 1196
rect 1194 1384 1206 1386
rect 1194 1376 1196 1384
rect 1204 1376 1206 1384
rect 874 1176 876 1184
rect 884 1176 886 1184
rect 874 1174 886 1176
rect 938 1184 950 1186
rect 938 1176 940 1184
rect 948 1176 950 1184
rect 810 1076 812 1084
rect 820 1076 822 1084
rect 810 1074 822 1076
rect 938 964 950 1176
rect 1194 1144 1206 1376
rect 1290 1204 1302 1456
rect 1450 1344 1462 1496
rect 1450 1336 1452 1344
rect 1460 1336 1462 1344
rect 1450 1334 1462 1336
rect 1290 1196 1292 1204
rect 1300 1196 1302 1204
rect 1290 1194 1302 1196
rect 1386 1304 1398 1306
rect 1386 1296 1388 1304
rect 1396 1296 1398 1304
rect 1194 1136 1196 1144
rect 1204 1136 1206 1144
rect 1194 1134 1206 1136
rect 938 956 940 964
rect 948 956 950 964
rect 938 954 950 956
rect 1066 984 1078 986
rect 1066 976 1068 984
rect 1076 976 1078 984
rect 650 496 652 504
rect 660 496 662 504
rect 650 494 662 496
rect 554 276 556 284
rect 564 276 566 284
rect 554 274 566 276
rect 1066 284 1078 976
rect 1322 904 1334 906
rect 1322 896 1324 904
rect 1332 896 1334 904
rect 1322 724 1334 896
rect 1386 864 1398 1296
rect 1560 1214 1608 1606
rect 1642 1984 1654 1986
rect 1642 1976 1644 1984
rect 1652 1976 1654 1984
rect 1642 1364 1654 1976
rect 1674 1784 1686 2356
rect 1674 1776 1676 1784
rect 1684 1776 1686 1784
rect 1674 1774 1686 1776
rect 1866 1724 1878 3356
rect 2826 3364 2838 3366
rect 2826 3356 2828 3364
rect 2836 3356 2838 3364
rect 2826 3284 2838 3356
rect 2826 3276 2828 3284
rect 2836 3276 2838 3284
rect 2826 3274 2838 3276
rect 1962 3264 1974 3266
rect 1962 3256 1964 3264
rect 1972 3256 1974 3264
rect 1930 3204 1942 3206
rect 1930 3196 1932 3204
rect 1940 3196 1942 3204
rect 1930 2664 1942 3196
rect 1962 2724 1974 3256
rect 1962 2716 1964 2724
rect 1972 2716 1974 2724
rect 1962 2714 1974 2716
rect 1994 3164 2006 3166
rect 1994 3156 1996 3164
rect 2004 3156 2006 3164
rect 1930 2656 1932 2664
rect 1940 2656 1942 2664
rect 1930 1784 1942 2656
rect 1994 2424 2006 3156
rect 2858 3084 2870 3636
rect 2922 3604 2934 3606
rect 2922 3596 2924 3604
rect 2932 3596 2934 3604
rect 2858 3076 2860 3084
rect 2868 3076 2870 3084
rect 2858 3074 2870 3076
rect 2890 3464 2902 3466
rect 2890 3456 2892 3464
rect 2900 3456 2902 3464
rect 2890 3064 2902 3456
rect 2922 3444 2934 3596
rect 2922 3436 2924 3444
rect 2932 3436 2934 3444
rect 2922 3434 2934 3436
rect 2954 3544 2966 3546
rect 2954 3536 2956 3544
rect 2964 3536 2966 3544
rect 2954 3444 2966 3536
rect 2954 3436 2956 3444
rect 2964 3436 2966 3444
rect 2954 3434 2966 3436
rect 3018 3484 3030 3486
rect 3018 3476 3020 3484
rect 3028 3476 3030 3484
rect 3018 3124 3030 3476
rect 3050 3364 3062 3716
rect 3082 3704 3094 3796
rect 3082 3696 3084 3704
rect 3092 3696 3094 3704
rect 3082 3694 3094 3696
rect 3050 3356 3052 3364
rect 3060 3356 3062 3364
rect 3050 3354 3062 3356
rect 3112 3414 3160 3806
rect 3112 3406 3116 3414
rect 3124 3406 3132 3414
rect 3140 3406 3148 3414
rect 3156 3406 3160 3414
rect 3018 3116 3020 3124
rect 3028 3116 3030 3124
rect 3018 3114 3030 3116
rect 2890 3056 2892 3064
rect 2900 3056 2902 3064
rect 2890 3054 2902 3056
rect 2922 3044 2934 3046
rect 2922 3036 2924 3044
rect 2932 3036 2934 3044
rect 2794 3024 2806 3026
rect 2794 3016 2796 3024
rect 2804 3016 2806 3024
rect 2698 2904 2710 2906
rect 2698 2896 2700 2904
rect 2708 2896 2710 2904
rect 1994 2416 1996 2424
rect 2004 2416 2006 2424
rect 1994 2414 2006 2416
rect 2058 2684 2070 2686
rect 2058 2676 2060 2684
rect 2068 2676 2070 2684
rect 2058 2284 2070 2676
rect 2506 2544 2518 2546
rect 2506 2536 2508 2544
rect 2516 2536 2518 2544
rect 2058 2276 2060 2284
rect 2068 2276 2070 2284
rect 2058 2274 2070 2276
rect 2250 2424 2262 2426
rect 2250 2416 2252 2424
rect 2260 2416 2262 2424
rect 2250 2184 2262 2416
rect 2506 2364 2518 2536
rect 2634 2444 2646 2446
rect 2634 2436 2636 2444
rect 2644 2436 2646 2444
rect 2506 2356 2508 2364
rect 2516 2356 2518 2364
rect 2506 2204 2518 2356
rect 2602 2424 2614 2426
rect 2602 2416 2604 2424
rect 2612 2416 2614 2424
rect 2602 2264 2614 2416
rect 2634 2344 2646 2436
rect 2698 2384 2710 2896
rect 2794 2824 2806 3016
rect 2794 2816 2796 2824
rect 2804 2816 2806 2824
rect 2794 2814 2806 2816
rect 2858 2964 2870 2966
rect 2858 2956 2860 2964
rect 2868 2956 2870 2964
rect 2762 2804 2774 2806
rect 2762 2796 2764 2804
rect 2772 2796 2774 2804
rect 2730 2684 2742 2686
rect 2730 2676 2732 2684
rect 2740 2676 2742 2684
rect 2730 2644 2742 2676
rect 2730 2636 2732 2644
rect 2740 2636 2742 2644
rect 2730 2634 2742 2636
rect 2698 2376 2700 2384
rect 2708 2376 2710 2384
rect 2698 2374 2710 2376
rect 2634 2336 2636 2344
rect 2644 2336 2646 2344
rect 2634 2334 2646 2336
rect 2666 2344 2678 2346
rect 2666 2336 2668 2344
rect 2676 2336 2678 2344
rect 2602 2256 2604 2264
rect 2612 2256 2614 2264
rect 2602 2254 2614 2256
rect 2506 2196 2508 2204
rect 2516 2196 2518 2204
rect 2506 2194 2518 2196
rect 2250 2176 2252 2184
rect 2260 2176 2262 2184
rect 2250 2174 2262 2176
rect 2346 2144 2358 2146
rect 2346 2136 2348 2144
rect 2356 2136 2358 2144
rect 2314 2104 2326 2106
rect 2314 2096 2316 2104
rect 2324 2096 2326 2104
rect 1930 1776 1932 1784
rect 1940 1776 1942 1784
rect 1930 1744 1942 1776
rect 1930 1736 1932 1744
rect 1940 1736 1942 1744
rect 1930 1734 1942 1736
rect 2058 1944 2070 1946
rect 2058 1936 2060 1944
rect 2068 1936 2070 1944
rect 2058 1744 2070 1936
rect 2058 1736 2060 1744
rect 2068 1736 2070 1744
rect 2058 1734 2070 1736
rect 2122 1924 2134 1926
rect 2122 1916 2124 1924
rect 2132 1916 2134 1924
rect 1866 1716 1868 1724
rect 1876 1716 1878 1724
rect 1866 1714 1878 1716
rect 1994 1644 2006 1646
rect 1994 1636 1996 1644
rect 2004 1636 2006 1644
rect 1642 1356 1644 1364
rect 1652 1356 1654 1364
rect 1642 1284 1654 1356
rect 1834 1424 1846 1426
rect 1834 1416 1836 1424
rect 1844 1416 1846 1424
rect 1642 1276 1644 1284
rect 1652 1276 1654 1284
rect 1642 1274 1654 1276
rect 1706 1284 1718 1286
rect 1706 1276 1708 1284
rect 1716 1276 1718 1284
rect 1560 1206 1564 1214
rect 1572 1206 1580 1214
rect 1588 1206 1596 1214
rect 1604 1206 1608 1214
rect 1386 856 1388 864
rect 1396 856 1398 864
rect 1386 854 1398 856
rect 1482 1064 1494 1066
rect 1482 1056 1484 1064
rect 1492 1056 1494 1064
rect 1322 716 1324 724
rect 1332 716 1334 724
rect 1322 714 1334 716
rect 1482 644 1494 1056
rect 1482 636 1484 644
rect 1492 636 1494 644
rect 1482 634 1494 636
rect 1560 814 1608 1206
rect 1706 1124 1718 1276
rect 1706 1116 1708 1124
rect 1716 1116 1718 1124
rect 1706 1114 1718 1116
rect 1834 1064 1846 1416
rect 1994 1264 2006 1636
rect 1994 1256 1996 1264
rect 2004 1256 2006 1264
rect 1994 1254 2006 1256
rect 2090 1364 2102 1366
rect 2090 1356 2092 1364
rect 2100 1356 2102 1364
rect 1930 1244 1942 1246
rect 1930 1236 1932 1244
rect 1940 1236 1942 1244
rect 1930 1184 1942 1236
rect 2090 1224 2102 1356
rect 2090 1216 2092 1224
rect 2100 1216 2102 1224
rect 2090 1214 2102 1216
rect 1930 1176 1932 1184
rect 1940 1176 1942 1184
rect 1930 1144 1942 1176
rect 1930 1136 1932 1144
rect 1940 1136 1942 1144
rect 1930 1134 1942 1136
rect 2122 1084 2134 1916
rect 2122 1076 2124 1084
rect 2132 1076 2134 1084
rect 2122 1074 2134 1076
rect 2154 1484 2166 1486
rect 2154 1476 2156 1484
rect 2164 1476 2166 1484
rect 1834 1056 1836 1064
rect 1844 1056 1846 1064
rect 1834 1054 1846 1056
rect 2154 924 2166 1476
rect 2250 1244 2262 1246
rect 2250 1236 2252 1244
rect 2260 1236 2262 1244
rect 2250 1024 2262 1236
rect 2250 1016 2252 1024
rect 2260 1016 2262 1024
rect 2250 1014 2262 1016
rect 2154 916 2156 924
rect 2164 916 2166 924
rect 2154 914 2166 916
rect 2314 924 2326 2096
rect 2346 1944 2358 2136
rect 2474 2064 2486 2066
rect 2474 2056 2476 2064
rect 2484 2056 2486 2064
rect 2346 1936 2348 1944
rect 2356 1936 2358 1944
rect 2346 1934 2358 1936
rect 2410 2004 2422 2006
rect 2410 1996 2412 2004
rect 2420 1996 2422 2004
rect 2346 1904 2358 1906
rect 2346 1896 2348 1904
rect 2356 1896 2358 1904
rect 2346 1864 2358 1896
rect 2346 1856 2348 1864
rect 2356 1856 2358 1864
rect 2346 1854 2358 1856
rect 2378 1844 2390 1846
rect 2378 1836 2380 1844
rect 2388 1836 2390 1844
rect 2346 1764 2358 1766
rect 2346 1756 2348 1764
rect 2356 1756 2358 1764
rect 2346 1524 2358 1756
rect 2346 1516 2348 1524
rect 2356 1516 2358 1524
rect 2346 1514 2358 1516
rect 2314 916 2316 924
rect 2324 916 2326 924
rect 2314 914 2326 916
rect 2346 1084 2358 1086
rect 2346 1076 2348 1084
rect 2356 1076 2358 1084
rect 1560 806 1564 814
rect 1572 806 1580 814
rect 1588 806 1596 814
rect 1604 806 1608 814
rect 1354 604 1366 606
rect 1354 596 1356 604
rect 1364 596 1366 604
rect 1322 584 1334 586
rect 1322 576 1324 584
rect 1332 576 1334 584
rect 1322 324 1334 576
rect 1322 316 1324 324
rect 1332 316 1334 324
rect 1322 314 1334 316
rect 1066 276 1068 284
rect 1076 276 1078 284
rect 1066 274 1078 276
rect 810 244 822 246
rect 810 236 812 244
rect 820 236 822 244
rect 714 164 726 166
rect 714 156 716 164
rect 724 156 726 164
rect 714 104 726 156
rect 810 144 822 236
rect 1354 244 1366 596
rect 1450 584 1462 586
rect 1450 576 1452 584
rect 1460 576 1462 584
rect 1450 444 1462 576
rect 1450 436 1452 444
rect 1460 436 1462 444
rect 1450 434 1462 436
rect 1354 236 1356 244
rect 1364 236 1366 244
rect 1354 234 1366 236
rect 1560 414 1608 806
rect 2346 804 2358 1076
rect 2378 904 2390 1836
rect 2378 896 2380 904
rect 2388 896 2390 904
rect 2378 894 2390 896
rect 2410 924 2422 1996
rect 2442 1944 2454 1946
rect 2442 1936 2444 1944
rect 2452 1936 2454 1944
rect 2442 1864 2454 1936
rect 2442 1856 2444 1864
rect 2452 1856 2454 1864
rect 2442 1854 2454 1856
rect 2474 1784 2486 2056
rect 2602 2064 2614 2066
rect 2602 2056 2604 2064
rect 2612 2056 2614 2064
rect 2474 1776 2476 1784
rect 2484 1776 2486 1784
rect 2474 1774 2486 1776
rect 2506 1804 2518 1806
rect 2506 1796 2508 1804
rect 2516 1796 2518 1804
rect 2442 1584 2454 1586
rect 2442 1576 2444 1584
rect 2452 1576 2454 1584
rect 2442 1324 2454 1576
rect 2506 1464 2518 1796
rect 2602 1764 2614 2056
rect 2602 1756 2604 1764
rect 2612 1756 2614 1764
rect 2602 1754 2614 1756
rect 2602 1704 2614 1706
rect 2602 1696 2604 1704
rect 2612 1696 2614 1704
rect 2602 1524 2614 1696
rect 2602 1516 2604 1524
rect 2612 1516 2614 1524
rect 2602 1514 2614 1516
rect 2666 1484 2678 2336
rect 2762 1944 2774 2796
rect 2826 2744 2838 2746
rect 2826 2736 2828 2744
rect 2836 2736 2838 2744
rect 2762 1936 2764 1944
rect 2772 1936 2774 1944
rect 2762 1934 2774 1936
rect 2794 2664 2806 2666
rect 2794 2656 2796 2664
rect 2804 2656 2806 2664
rect 2794 1784 2806 2656
rect 2826 2524 2838 2736
rect 2858 2724 2870 2956
rect 2858 2716 2860 2724
rect 2868 2716 2870 2724
rect 2858 2714 2870 2716
rect 2826 2516 2828 2524
rect 2836 2516 2838 2524
rect 2826 2514 2838 2516
rect 2922 2504 2934 3036
rect 3112 3014 3160 3406
rect 3112 3006 3116 3014
rect 3124 3006 3132 3014
rect 3140 3006 3148 3014
rect 3156 3006 3160 3014
rect 2954 2964 2966 2966
rect 2954 2956 2956 2964
rect 2964 2956 2966 2964
rect 2954 2804 2966 2956
rect 2954 2796 2956 2804
rect 2964 2796 2966 2804
rect 2954 2794 2966 2796
rect 3082 2804 3094 2806
rect 3082 2796 3084 2804
rect 3092 2796 3094 2804
rect 2986 2644 2998 2646
rect 2986 2636 2988 2644
rect 2996 2636 2998 2644
rect 2922 2496 2924 2504
rect 2932 2496 2934 2504
rect 2922 2494 2934 2496
rect 2954 2504 2966 2506
rect 2954 2496 2956 2504
rect 2964 2496 2966 2504
rect 2858 2484 2870 2486
rect 2858 2476 2860 2484
rect 2868 2476 2870 2484
rect 2858 2304 2870 2476
rect 2954 2424 2966 2496
rect 2954 2416 2956 2424
rect 2964 2416 2966 2424
rect 2954 2414 2966 2416
rect 2986 2424 2998 2636
rect 2986 2416 2988 2424
rect 2996 2416 2998 2424
rect 2986 2414 2998 2416
rect 3050 2404 3062 2406
rect 3050 2396 3052 2404
rect 3060 2396 3062 2404
rect 2858 2296 2860 2304
rect 2868 2296 2870 2304
rect 2858 2294 2870 2296
rect 3018 2324 3030 2326
rect 3018 2316 3020 2324
rect 3028 2316 3030 2324
rect 3018 2284 3030 2316
rect 3018 2276 3020 2284
rect 3028 2276 3030 2284
rect 3018 2274 3030 2276
rect 2922 2224 2934 2226
rect 2922 2216 2924 2224
rect 2932 2216 2934 2224
rect 2890 2204 2902 2206
rect 2890 2196 2892 2204
rect 2900 2196 2902 2204
rect 2794 1776 2796 1784
rect 2804 1776 2806 1784
rect 2794 1774 2806 1776
rect 2826 2124 2838 2126
rect 2826 2116 2828 2124
rect 2836 2116 2838 2124
rect 2666 1476 2668 1484
rect 2676 1476 2678 1484
rect 2666 1474 2678 1476
rect 2794 1564 2806 1566
rect 2794 1556 2796 1564
rect 2804 1556 2806 1564
rect 2506 1456 2508 1464
rect 2516 1456 2518 1464
rect 2506 1454 2518 1456
rect 2794 1404 2806 1556
rect 2794 1396 2796 1404
rect 2804 1396 2806 1404
rect 2794 1394 2806 1396
rect 2442 1316 2444 1324
rect 2452 1316 2454 1324
rect 2442 1314 2454 1316
rect 2666 1364 2678 1366
rect 2666 1356 2668 1364
rect 2676 1356 2678 1364
rect 2410 916 2412 924
rect 2420 916 2422 924
rect 2346 796 2348 804
rect 2356 796 2358 804
rect 2346 794 2358 796
rect 2410 664 2422 916
rect 2442 1124 2454 1126
rect 2442 1116 2444 1124
rect 2452 1116 2454 1124
rect 2442 844 2454 1116
rect 2442 836 2444 844
rect 2452 836 2454 844
rect 2442 834 2454 836
rect 2474 1044 2486 1046
rect 2474 1036 2476 1044
rect 2484 1036 2486 1044
rect 2410 656 2412 664
rect 2420 656 2422 664
rect 2410 654 2422 656
rect 2474 664 2486 1036
rect 2474 656 2476 664
rect 2484 656 2486 664
rect 2474 654 2486 656
rect 2506 1004 2518 1006
rect 2506 996 2508 1004
rect 2516 996 2518 1004
rect 2506 604 2518 996
rect 2666 944 2678 1356
rect 2666 936 2668 944
rect 2676 936 2678 944
rect 2666 934 2678 936
rect 2730 1304 2742 1306
rect 2730 1296 2732 1304
rect 2740 1296 2742 1304
rect 2506 596 2508 604
rect 2516 596 2518 604
rect 2506 594 2518 596
rect 2602 924 2614 926
rect 2602 916 2604 924
rect 2612 916 2614 924
rect 1560 406 1564 414
rect 1572 406 1580 414
rect 1588 406 1596 414
rect 1604 406 1608 414
rect 810 136 812 144
rect 820 136 822 144
rect 810 134 822 136
rect 714 96 716 104
rect 724 96 726 104
rect 714 94 726 96
rect 1560 14 1608 406
rect 2154 264 2166 266
rect 2154 256 2156 264
rect 2164 256 2166 264
rect 1930 124 2038 126
rect 1930 116 2028 124
rect 2036 116 2038 124
rect 1930 114 2038 116
rect 1930 104 1942 114
rect 1930 96 1932 104
rect 1940 96 1942 104
rect 1930 94 1942 96
rect 2154 24 2166 256
rect 2154 16 2156 24
rect 2164 16 2166 24
rect 2154 14 2166 16
rect 2314 264 2326 266
rect 2314 256 2316 264
rect 2324 256 2326 264
rect 2314 24 2326 256
rect 2314 16 2316 24
rect 2324 16 2326 24
rect 2314 14 2326 16
rect 2602 24 2614 916
rect 2730 804 2742 1296
rect 2762 1264 2774 1266
rect 2762 1256 2764 1264
rect 2772 1256 2774 1264
rect 2762 1024 2774 1256
rect 2762 1016 2764 1024
rect 2772 1016 2774 1024
rect 2762 1014 2774 1016
rect 2826 964 2838 2116
rect 2826 956 2828 964
rect 2836 956 2838 964
rect 2826 954 2838 956
rect 2858 2064 2870 2066
rect 2858 2056 2860 2064
rect 2868 2056 2870 2064
rect 2858 904 2870 2056
rect 2858 896 2860 904
rect 2868 896 2870 904
rect 2858 894 2870 896
rect 2890 904 2902 2196
rect 2922 1964 2934 2216
rect 3050 2164 3062 2396
rect 3050 2156 3052 2164
rect 3060 2156 3062 2164
rect 3050 2154 3062 2156
rect 3018 2144 3030 2146
rect 3018 2136 3020 2144
rect 3028 2136 3030 2144
rect 2922 1956 2924 1964
rect 2932 1956 2934 1964
rect 2922 1954 2934 1956
rect 2954 2084 2966 2086
rect 2954 2076 2956 2084
rect 2964 2076 2966 2084
rect 2954 1864 2966 2076
rect 3018 2044 3030 2136
rect 3018 2036 3020 2044
rect 3028 2036 3030 2044
rect 3018 2034 3030 2036
rect 2954 1856 2956 1864
rect 2964 1856 2966 1864
rect 2954 1854 2966 1856
rect 3050 1984 3062 1986
rect 3050 1976 3052 1984
rect 3060 1976 3062 1984
rect 3018 1744 3030 1746
rect 3018 1736 3020 1744
rect 3028 1736 3030 1744
rect 3018 1664 3030 1736
rect 3050 1744 3062 1976
rect 3082 1804 3094 2796
rect 3082 1796 3084 1804
rect 3092 1796 3094 1804
rect 3082 1794 3094 1796
rect 3112 2614 3160 3006
rect 3112 2606 3116 2614
rect 3124 2606 3132 2614
rect 3140 2606 3148 2614
rect 3156 2606 3160 2614
rect 3112 2214 3160 2606
rect 3178 3844 3190 3846
rect 3178 3836 3180 3844
rect 3188 3836 3190 3844
rect 3178 2564 3190 3836
rect 3210 3204 3222 3856
rect 3274 3844 3286 4156
rect 3274 3836 3276 3844
rect 3284 3836 3286 3844
rect 3274 3834 3286 3836
rect 3338 4104 3350 4106
rect 3338 4096 3340 4104
rect 3348 4096 3350 4104
rect 3306 3784 3318 3786
rect 3306 3776 3308 3784
rect 3316 3776 3318 3784
rect 3210 3196 3212 3204
rect 3220 3196 3222 3204
rect 3210 3194 3222 3196
rect 3274 3604 3286 3606
rect 3274 3596 3276 3604
rect 3284 3596 3286 3604
rect 3274 3144 3286 3596
rect 3274 3136 3276 3144
rect 3284 3136 3286 3144
rect 3274 3134 3286 3136
rect 3242 3124 3254 3126
rect 3242 3116 3244 3124
rect 3252 3116 3254 3124
rect 3178 2556 3180 2564
rect 3188 2556 3190 2564
rect 3178 2554 3190 2556
rect 3210 3044 3222 3046
rect 3210 3036 3212 3044
rect 3220 3036 3222 3044
rect 3210 2684 3222 3036
rect 3210 2676 3212 2684
rect 3220 2676 3222 2684
rect 3112 2206 3116 2214
rect 3124 2206 3132 2214
rect 3140 2206 3148 2214
rect 3156 2206 3160 2214
rect 3112 1814 3160 2206
rect 3178 2304 3190 2306
rect 3178 2296 3180 2304
rect 3188 2296 3190 2304
rect 3178 2064 3190 2296
rect 3178 2056 3180 2064
rect 3188 2056 3190 2064
rect 3178 2024 3190 2056
rect 3178 2016 3180 2024
rect 3188 2016 3190 2024
rect 3178 2014 3190 2016
rect 3112 1806 3116 1814
rect 3124 1806 3132 1814
rect 3140 1806 3148 1814
rect 3156 1806 3160 1814
rect 3050 1736 3052 1744
rect 3060 1736 3062 1744
rect 3050 1734 3062 1736
rect 3082 1764 3094 1766
rect 3082 1756 3084 1764
rect 3092 1756 3094 1764
rect 3018 1656 3020 1664
rect 3028 1656 3030 1664
rect 3018 1654 3030 1656
rect 2986 1564 2998 1566
rect 2986 1556 2988 1564
rect 2996 1556 2998 1564
rect 2954 1544 2966 1546
rect 2954 1536 2956 1544
rect 2964 1536 2966 1544
rect 2954 1424 2966 1536
rect 2954 1416 2956 1424
rect 2964 1416 2966 1424
rect 2954 1414 2966 1416
rect 2986 1424 2998 1556
rect 2986 1416 2988 1424
rect 2996 1416 2998 1424
rect 2986 1414 2998 1416
rect 3050 1424 3062 1426
rect 3050 1416 3052 1424
rect 3060 1416 3062 1424
rect 2954 1344 2966 1346
rect 2954 1336 2956 1344
rect 2964 1336 2966 1344
rect 2890 896 2892 904
rect 2900 896 2902 904
rect 2890 894 2902 896
rect 2922 1224 2934 1226
rect 2922 1216 2924 1224
rect 2932 1216 2934 1224
rect 2922 884 2934 1216
rect 2922 876 2924 884
rect 2932 876 2934 884
rect 2922 874 2934 876
rect 2954 824 2966 1336
rect 3018 1304 3030 1306
rect 3018 1296 3020 1304
rect 3028 1296 3030 1304
rect 2986 1004 2998 1006
rect 2986 996 2988 1004
rect 2996 996 2998 1004
rect 2986 964 2998 996
rect 2986 956 2988 964
rect 2996 956 2998 964
rect 2986 954 2998 956
rect 3018 844 3030 1296
rect 3018 836 3020 844
rect 3028 836 3030 844
rect 3018 834 3030 836
rect 2954 816 2956 824
rect 2964 816 2966 824
rect 2954 814 2966 816
rect 2986 824 2998 826
rect 2986 816 2988 824
rect 2996 816 2998 824
rect 2730 796 2732 804
rect 2740 796 2742 804
rect 2730 794 2742 796
rect 2698 724 2710 726
rect 2698 716 2700 724
rect 2708 716 2710 724
rect 2698 64 2710 716
rect 2986 624 2998 816
rect 3050 824 3062 1416
rect 3082 1364 3094 1756
rect 3082 1356 3084 1364
rect 3092 1356 3094 1364
rect 3082 1354 3094 1356
rect 3112 1414 3160 1806
rect 3178 1864 3190 1866
rect 3178 1856 3180 1864
rect 3188 1856 3190 1864
rect 3178 1804 3190 1856
rect 3178 1796 3180 1804
rect 3188 1796 3190 1804
rect 3178 1794 3190 1796
rect 3112 1406 3116 1414
rect 3124 1406 3132 1414
rect 3140 1406 3148 1414
rect 3156 1406 3160 1414
rect 3050 816 3052 824
rect 3060 816 3062 824
rect 3050 814 3062 816
rect 3112 1014 3160 1406
rect 3112 1006 3116 1014
rect 3124 1006 3132 1014
rect 3140 1006 3148 1014
rect 3156 1006 3160 1014
rect 2986 616 2988 624
rect 2996 616 2998 624
rect 2986 614 2998 616
rect 3112 614 3160 1006
rect 3178 1744 3190 1746
rect 3178 1736 3180 1744
rect 3188 1736 3190 1744
rect 3178 1504 3190 1736
rect 3210 1744 3222 2676
rect 3242 2404 3254 3116
rect 3274 3064 3286 3066
rect 3274 3056 3276 3064
rect 3284 3056 3286 3064
rect 3274 2884 3286 3056
rect 3274 2876 3276 2884
rect 3284 2876 3286 2884
rect 3274 2874 3286 2876
rect 3242 2396 3244 2404
rect 3252 2396 3254 2404
rect 3242 2394 3254 2396
rect 3306 2524 3318 3776
rect 3338 3764 3350 4096
rect 3370 4084 3382 4376
rect 3402 4364 3414 4936
rect 3434 4704 3446 4706
rect 3434 4696 3436 4704
rect 3444 4696 3446 4704
rect 3434 4464 3446 4696
rect 3434 4456 3436 4464
rect 3444 4456 3446 4464
rect 3434 4454 3446 4456
rect 3402 4356 3404 4364
rect 3412 4356 3414 4364
rect 3402 4354 3414 4356
rect 3370 4076 3372 4084
rect 3380 4076 3382 4084
rect 3370 4074 3382 4076
rect 3434 4344 3446 4346
rect 3434 4336 3436 4344
rect 3444 4336 3446 4344
rect 3434 3904 3446 4336
rect 3466 4044 3478 5116
rect 3498 5044 3510 5336
rect 3562 5184 3574 5376
rect 3690 5324 3702 5326
rect 3690 5316 3692 5324
rect 3700 5316 3702 5324
rect 3690 5284 3702 5316
rect 3690 5276 3692 5284
rect 3700 5276 3702 5284
rect 3690 5274 3702 5276
rect 3562 5176 3564 5184
rect 3572 5176 3574 5184
rect 3562 5086 3574 5176
rect 3562 5084 3590 5086
rect 3562 5076 3580 5084
rect 3588 5076 3590 5084
rect 3562 5074 3590 5076
rect 3498 5036 3500 5044
rect 3508 5036 3510 5044
rect 3498 5034 3510 5036
rect 3530 4884 3542 4886
rect 3530 4876 3532 4884
rect 3540 4876 3542 4884
rect 3530 4484 3542 4876
rect 3530 4476 3532 4484
rect 3540 4476 3542 4484
rect 3530 4474 3542 4476
rect 3594 4504 3606 4506
rect 3594 4496 3596 4504
rect 3604 4496 3606 4504
rect 3466 4036 3468 4044
rect 3476 4036 3478 4044
rect 3466 4034 3478 4036
rect 3562 4264 3574 4266
rect 3562 4256 3564 4264
rect 3572 4256 3574 4264
rect 3434 3896 3436 3904
rect 3444 3896 3446 3904
rect 3434 3894 3446 3896
rect 3562 3864 3574 4256
rect 3562 3856 3564 3864
rect 3572 3856 3574 3864
rect 3562 3854 3574 3856
rect 3594 4064 3606 4496
rect 3594 4056 3596 4064
rect 3604 4056 3606 4064
rect 3338 3756 3340 3764
rect 3348 3756 3350 3764
rect 3338 3624 3350 3756
rect 3498 3824 3510 3826
rect 3498 3816 3500 3824
rect 3508 3816 3510 3824
rect 3498 3684 3510 3816
rect 3498 3676 3500 3684
rect 3508 3676 3510 3684
rect 3498 3674 3510 3676
rect 3562 3784 3574 3786
rect 3562 3776 3564 3784
rect 3572 3776 3574 3784
rect 3338 3616 3340 3624
rect 3348 3616 3350 3624
rect 3338 3124 3350 3616
rect 3530 3504 3542 3506
rect 3530 3496 3532 3504
rect 3540 3496 3542 3504
rect 3402 3484 3414 3486
rect 3402 3476 3404 3484
rect 3412 3476 3414 3484
rect 3402 3324 3414 3476
rect 3498 3484 3510 3486
rect 3498 3476 3500 3484
rect 3508 3476 3510 3484
rect 3402 3316 3404 3324
rect 3412 3316 3414 3324
rect 3402 3314 3414 3316
rect 3434 3384 3446 3386
rect 3434 3376 3436 3384
rect 3444 3376 3446 3384
rect 3338 3116 3340 3124
rect 3348 3116 3350 3124
rect 3338 3114 3350 3116
rect 3370 3304 3382 3306
rect 3370 3296 3372 3304
rect 3380 3296 3382 3304
rect 3370 2924 3382 3296
rect 3434 3164 3446 3376
rect 3498 3224 3510 3476
rect 3530 3324 3542 3496
rect 3562 3364 3574 3776
rect 3594 3784 3606 4056
rect 3594 3776 3596 3784
rect 3604 3776 3606 3784
rect 3594 3774 3606 3776
rect 3626 4264 3638 4266
rect 3626 4256 3628 4264
rect 3636 4256 3638 4264
rect 3562 3356 3564 3364
rect 3572 3356 3574 3364
rect 3562 3354 3574 3356
rect 3594 3724 3606 3726
rect 3594 3716 3596 3724
rect 3604 3716 3606 3724
rect 3530 3316 3532 3324
rect 3540 3316 3542 3324
rect 3530 3314 3542 3316
rect 3498 3216 3500 3224
rect 3508 3216 3510 3224
rect 3498 3214 3510 3216
rect 3434 3156 3436 3164
rect 3444 3156 3446 3164
rect 3434 3154 3446 3156
rect 3370 2916 3372 2924
rect 3380 2916 3382 2924
rect 3370 2914 3382 2916
rect 3562 3084 3574 3086
rect 3562 3076 3564 3084
rect 3572 3076 3574 3084
rect 3562 2944 3574 3076
rect 3562 2936 3564 2944
rect 3572 2936 3574 2944
rect 3370 2844 3382 2846
rect 3370 2836 3372 2844
rect 3380 2836 3382 2844
rect 3370 2784 3382 2836
rect 3370 2776 3372 2784
rect 3380 2776 3382 2784
rect 3370 2774 3382 2776
rect 3466 2824 3478 2826
rect 3466 2816 3468 2824
rect 3476 2816 3478 2824
rect 3402 2744 3414 2746
rect 3402 2736 3404 2744
rect 3412 2736 3414 2744
rect 3306 2516 3308 2524
rect 3316 2516 3318 2524
rect 3274 2364 3286 2366
rect 3274 2356 3276 2364
rect 3284 2356 3286 2364
rect 3242 2304 3254 2306
rect 3242 2296 3244 2304
rect 3252 2296 3254 2304
rect 3242 2124 3254 2296
rect 3242 2116 3244 2124
rect 3252 2116 3254 2124
rect 3242 2114 3254 2116
rect 3274 1884 3286 2356
rect 3274 1876 3276 1884
rect 3284 1876 3286 1884
rect 3274 1874 3286 1876
rect 3306 2284 3318 2516
rect 3338 2624 3350 2626
rect 3338 2616 3340 2624
rect 3348 2616 3350 2624
rect 3338 2404 3350 2616
rect 3370 2544 3382 2546
rect 3370 2536 3372 2544
rect 3380 2536 3382 2544
rect 3370 2464 3382 2536
rect 3402 2544 3414 2736
rect 3466 2724 3478 2816
rect 3466 2716 3468 2724
rect 3476 2716 3478 2724
rect 3466 2714 3478 2716
rect 3498 2824 3510 2826
rect 3498 2816 3500 2824
rect 3508 2816 3510 2824
rect 3402 2536 3404 2544
rect 3412 2536 3414 2544
rect 3402 2534 3414 2536
rect 3466 2684 3478 2686
rect 3466 2676 3468 2684
rect 3476 2676 3478 2684
rect 3466 2484 3478 2676
rect 3498 2664 3510 2816
rect 3498 2656 3500 2664
rect 3508 2656 3510 2664
rect 3498 2654 3510 2656
rect 3466 2476 3468 2484
rect 3476 2476 3478 2484
rect 3466 2474 3478 2476
rect 3530 2584 3542 2586
rect 3530 2576 3532 2584
rect 3540 2576 3542 2584
rect 3530 2484 3542 2576
rect 3530 2476 3532 2484
rect 3540 2476 3542 2484
rect 3530 2474 3542 2476
rect 3370 2456 3372 2464
rect 3380 2456 3382 2464
rect 3370 2454 3382 2456
rect 3338 2396 3340 2404
rect 3348 2396 3350 2404
rect 3338 2304 3350 2396
rect 3434 2424 3446 2426
rect 3434 2416 3436 2424
rect 3444 2416 3446 2424
rect 3338 2296 3340 2304
rect 3348 2296 3350 2304
rect 3338 2294 3350 2296
rect 3402 2304 3414 2306
rect 3402 2296 3404 2304
rect 3412 2296 3414 2304
rect 3306 2276 3308 2284
rect 3316 2276 3318 2284
rect 3210 1736 3212 1744
rect 3220 1736 3222 1744
rect 3210 1734 3222 1736
rect 3274 1784 3286 1786
rect 3274 1776 3276 1784
rect 3284 1776 3286 1784
rect 3178 1496 3180 1504
rect 3188 1496 3190 1504
rect 3178 1464 3190 1496
rect 3178 1456 3180 1464
rect 3188 1456 3190 1464
rect 3178 1344 3190 1456
rect 3178 1336 3180 1344
rect 3188 1336 3190 1344
rect 3178 924 3190 1336
rect 3210 1584 3222 1586
rect 3210 1576 3212 1584
rect 3220 1576 3222 1584
rect 3210 1344 3222 1576
rect 3274 1524 3286 1776
rect 3274 1516 3276 1524
rect 3284 1516 3286 1524
rect 3274 1484 3286 1516
rect 3274 1476 3276 1484
rect 3284 1476 3286 1484
rect 3274 1474 3286 1476
rect 3306 1784 3318 2276
rect 3370 2204 3382 2206
rect 3370 2196 3372 2204
rect 3380 2196 3382 2204
rect 3306 1776 3308 1784
rect 3316 1776 3318 1784
rect 3274 1424 3286 1426
rect 3274 1416 3276 1424
rect 3284 1416 3286 1424
rect 3210 1336 3212 1344
rect 3220 1336 3222 1344
rect 3210 1334 3222 1336
rect 3242 1344 3254 1346
rect 3242 1336 3244 1344
rect 3252 1336 3254 1344
rect 3178 916 3180 924
rect 3188 916 3190 924
rect 3178 914 3190 916
rect 3210 1164 3222 1166
rect 3210 1156 3212 1164
rect 3220 1156 3222 1164
rect 3210 884 3222 1156
rect 3242 1004 3254 1336
rect 3274 1164 3286 1416
rect 3274 1156 3276 1164
rect 3284 1156 3286 1164
rect 3274 1154 3286 1156
rect 3306 1064 3318 1776
rect 3338 2164 3350 2166
rect 3338 2156 3340 2164
rect 3348 2156 3350 2164
rect 3338 1264 3350 2156
rect 3370 2064 3382 2196
rect 3402 2084 3414 2296
rect 3402 2076 3404 2084
rect 3412 2076 3414 2084
rect 3402 2074 3414 2076
rect 3370 2056 3372 2064
rect 3380 2056 3382 2064
rect 3370 2054 3382 2056
rect 3402 1724 3414 1726
rect 3402 1716 3404 1724
rect 3412 1716 3414 1724
rect 3402 1384 3414 1716
rect 3434 1664 3446 2416
rect 3434 1656 3436 1664
rect 3444 1656 3446 1664
rect 3434 1654 3446 1656
rect 3466 2344 3478 2346
rect 3466 2336 3468 2344
rect 3476 2336 3478 2344
rect 3466 2164 3478 2336
rect 3466 2156 3468 2164
rect 3476 2156 3478 2164
rect 3466 1524 3478 2156
rect 3530 2324 3542 2326
rect 3530 2316 3532 2324
rect 3540 2316 3542 2324
rect 3498 2144 3510 2146
rect 3498 2136 3500 2144
rect 3508 2136 3510 2144
rect 3498 1784 3510 2136
rect 3530 2004 3542 2316
rect 3530 1996 3532 2004
rect 3540 1996 3542 2004
rect 3530 1994 3542 1996
rect 3562 2184 3574 2936
rect 3562 2176 3564 2184
rect 3572 2176 3574 2184
rect 3498 1776 3500 1784
rect 3508 1776 3510 1784
rect 3498 1774 3510 1776
rect 3562 1884 3574 2176
rect 3562 1876 3564 1884
rect 3572 1876 3574 1884
rect 3466 1516 3468 1524
rect 3476 1516 3478 1524
rect 3466 1514 3478 1516
rect 3402 1376 3404 1384
rect 3412 1376 3414 1384
rect 3402 1374 3414 1376
rect 3434 1504 3446 1506
rect 3434 1496 3436 1504
rect 3444 1496 3446 1504
rect 3338 1256 3340 1264
rect 3348 1256 3350 1264
rect 3338 1254 3350 1256
rect 3306 1056 3308 1064
rect 3316 1056 3318 1064
rect 3306 1054 3318 1056
rect 3242 996 3244 1004
rect 3252 996 3254 1004
rect 3242 994 3254 996
rect 3434 904 3446 1496
rect 3562 1484 3574 1876
rect 3594 3064 3606 3716
rect 3626 3384 3638 4256
rect 3658 4124 3670 4126
rect 3658 4116 3660 4124
rect 3668 4116 3670 4124
rect 3658 3744 3670 4116
rect 3658 3736 3660 3744
rect 3668 3736 3670 3744
rect 3658 3734 3670 3736
rect 3626 3376 3628 3384
rect 3636 3376 3638 3384
rect 3626 3374 3638 3376
rect 3690 3524 3702 3526
rect 3690 3516 3692 3524
rect 3700 3516 3702 3524
rect 3690 3384 3702 3516
rect 3722 3524 3734 5596
rect 3946 5484 3958 5486
rect 3946 5476 3948 5484
rect 3956 5476 3958 5484
rect 3754 5444 3766 5446
rect 3754 5436 3756 5444
rect 3764 5436 3766 5444
rect 3754 4664 3766 5436
rect 3946 5184 3958 5476
rect 4586 5344 4598 5346
rect 4586 5336 4588 5344
rect 4596 5336 4598 5344
rect 3946 5176 3948 5184
rect 3956 5176 3958 5184
rect 3946 5174 3958 5176
rect 4042 5244 4054 5246
rect 4042 5236 4044 5244
rect 4052 5236 4054 5244
rect 3882 5064 3894 5066
rect 3882 5056 3884 5064
rect 3892 5056 3894 5064
rect 3850 5044 3862 5046
rect 3850 5036 3852 5044
rect 3860 5036 3862 5044
rect 3850 4944 3862 5036
rect 3850 4936 3852 4944
rect 3860 4936 3862 4944
rect 3850 4934 3862 4936
rect 3850 4704 3862 4706
rect 3850 4696 3852 4704
rect 3860 4696 3862 4704
rect 3850 4686 3862 4696
rect 3754 4656 3756 4664
rect 3764 4656 3766 4664
rect 3754 4564 3766 4656
rect 3818 4674 3862 4686
rect 3818 4664 3830 4674
rect 3818 4656 3820 4664
rect 3828 4656 3830 4664
rect 3818 4654 3830 4656
rect 3882 4624 3894 5056
rect 4042 4924 4054 5236
rect 4362 5164 4374 5166
rect 4362 5156 4364 5164
rect 4372 5156 4374 5164
rect 4042 4916 4044 4924
rect 4052 4916 4054 4924
rect 4042 4914 4054 4916
rect 4202 4924 4214 4926
rect 4202 4916 4204 4924
rect 4212 4916 4214 4924
rect 3882 4616 3884 4624
rect 3892 4616 3894 4624
rect 3882 4614 3894 4616
rect 4042 4724 4054 4726
rect 4042 4716 4044 4724
rect 4052 4716 4054 4724
rect 3754 4556 3756 4564
rect 3764 4556 3766 4564
rect 3754 4554 3766 4556
rect 4042 4244 4054 4716
rect 4202 4444 4214 4916
rect 4202 4436 4204 4444
rect 4212 4436 4214 4444
rect 4202 4434 4214 4436
rect 4042 4236 4044 4244
rect 4052 4236 4054 4244
rect 4042 4234 4054 4236
rect 4234 4204 4246 4206
rect 4234 4196 4236 4204
rect 4244 4196 4246 4204
rect 3722 3516 3724 3524
rect 3732 3516 3734 3524
rect 3722 3514 3734 3516
rect 3754 4044 3766 4046
rect 3754 4036 3756 4044
rect 3764 4036 3766 4044
rect 3754 3404 3766 4036
rect 3850 3924 3862 3926
rect 3850 3916 3852 3924
rect 3860 3916 3862 3924
rect 3850 3804 3862 3916
rect 4234 3884 4246 4196
rect 4234 3876 4236 3884
rect 4244 3876 4246 3884
rect 4234 3874 4246 3876
rect 4266 4104 4278 4106
rect 4266 4096 4268 4104
rect 4276 4096 4278 4104
rect 4266 3884 4278 4096
rect 4266 3876 4268 3884
rect 4276 3876 4278 3884
rect 4266 3874 4278 3876
rect 4330 4104 4342 4106
rect 4330 4096 4332 4104
rect 4340 4096 4342 4104
rect 4330 3884 4342 4096
rect 4330 3876 4332 3884
rect 4340 3876 4342 3884
rect 4330 3874 4342 3876
rect 3850 3796 3852 3804
rect 3860 3796 3862 3804
rect 3850 3794 3862 3796
rect 4010 3844 4022 3846
rect 4010 3836 4012 3844
rect 4020 3836 4022 3844
rect 3754 3396 3756 3404
rect 3764 3396 3766 3404
rect 3754 3394 3766 3396
rect 3690 3376 3692 3384
rect 3700 3376 3702 3384
rect 3690 3374 3702 3376
rect 3658 3364 3670 3366
rect 3658 3356 3660 3364
rect 3668 3356 3670 3364
rect 3594 3056 3596 3064
rect 3604 3056 3606 3064
rect 3594 2604 3606 3056
rect 3626 3064 3638 3066
rect 3626 3056 3628 3064
rect 3636 3056 3638 3064
rect 3626 2744 3638 3056
rect 3626 2736 3628 2744
rect 3636 2736 3638 2744
rect 3626 2734 3638 2736
rect 3594 2596 3596 2604
rect 3604 2596 3606 2604
rect 3594 1864 3606 2596
rect 3626 2704 3638 2706
rect 3626 2696 3628 2704
rect 3636 2696 3638 2704
rect 3626 2544 3638 2696
rect 3626 2536 3628 2544
rect 3636 2536 3638 2544
rect 3626 2534 3638 2536
rect 3594 1856 3596 1864
rect 3604 1856 3606 1864
rect 3594 1854 3606 1856
rect 3658 1744 3670 3356
rect 3850 3304 3862 3306
rect 3850 3296 3852 3304
rect 3860 3296 3862 3304
rect 3754 3224 3766 3226
rect 3754 3216 3756 3224
rect 3764 3216 3766 3224
rect 3754 3084 3766 3216
rect 3754 3076 3756 3084
rect 3764 3076 3766 3084
rect 3754 3074 3766 3076
rect 3786 3104 3798 3106
rect 3786 3096 3788 3104
rect 3796 3096 3798 3104
rect 3786 3064 3798 3096
rect 3786 3056 3788 3064
rect 3796 3056 3798 3064
rect 3722 3044 3734 3046
rect 3722 3036 3724 3044
rect 3732 3036 3734 3044
rect 3722 2924 3734 3036
rect 3754 3024 3766 3026
rect 3754 3016 3756 3024
rect 3764 3016 3766 3024
rect 3754 2944 3766 3016
rect 3754 2936 3756 2944
rect 3764 2936 3766 2944
rect 3754 2934 3766 2936
rect 3722 2916 3724 2924
rect 3732 2916 3734 2924
rect 3722 2914 3734 2916
rect 3690 2864 3702 2866
rect 3690 2856 3692 2864
rect 3700 2856 3702 2864
rect 3690 2584 3702 2856
rect 3754 2864 3766 2866
rect 3754 2856 3756 2864
rect 3764 2856 3766 2864
rect 3754 2704 3766 2856
rect 3754 2696 3756 2704
rect 3764 2696 3766 2704
rect 3754 2694 3766 2696
rect 3786 2664 3798 3056
rect 3786 2656 3788 2664
rect 3796 2656 3798 2664
rect 3786 2654 3798 2656
rect 3690 2576 3692 2584
rect 3700 2576 3702 2584
rect 3690 2574 3702 2576
rect 3786 2624 3798 2626
rect 3786 2616 3788 2624
rect 3796 2616 3798 2624
rect 3786 2504 3798 2616
rect 3786 2496 3788 2504
rect 3796 2496 3798 2504
rect 3786 2494 3798 2496
rect 3850 2504 3862 3296
rect 4010 3044 4022 3836
rect 4202 3664 4214 3666
rect 4202 3656 4204 3664
rect 4212 3656 4214 3664
rect 4138 3564 4150 3566
rect 4138 3556 4140 3564
rect 4148 3556 4150 3564
rect 4138 3464 4150 3556
rect 4138 3456 4140 3464
rect 4148 3456 4150 3464
rect 4010 3036 4012 3044
rect 4020 3036 4022 3044
rect 4010 3034 4022 3036
rect 4074 3064 4086 3066
rect 4074 3056 4076 3064
rect 4084 3056 4086 3064
rect 3914 3004 3926 3006
rect 3914 2996 3916 3004
rect 3924 2996 3926 3004
rect 3914 2864 3926 2996
rect 3914 2856 3916 2864
rect 3924 2856 3926 2864
rect 3914 2854 3926 2856
rect 3882 2824 3894 2826
rect 3882 2816 3884 2824
rect 3892 2816 3894 2824
rect 3882 2664 3894 2816
rect 4042 2724 4054 2726
rect 4042 2716 4044 2724
rect 4052 2716 4054 2724
rect 3882 2656 3884 2664
rect 3892 2656 3894 2664
rect 3882 2654 3894 2656
rect 3914 2704 3926 2706
rect 3914 2696 3916 2704
rect 3924 2696 3926 2704
rect 3850 2496 3852 2504
rect 3860 2496 3862 2504
rect 3754 2424 3766 2426
rect 3754 2416 3756 2424
rect 3764 2416 3766 2424
rect 3754 2184 3766 2416
rect 3818 2424 3830 2426
rect 3818 2416 3820 2424
rect 3828 2416 3830 2424
rect 3818 2384 3830 2416
rect 3818 2376 3820 2384
rect 3828 2376 3830 2384
rect 3818 2374 3830 2376
rect 3754 2176 3756 2184
rect 3764 2176 3766 2184
rect 3754 2174 3766 2176
rect 3818 2004 3830 2006
rect 3818 1996 3820 2004
rect 3828 1996 3830 2004
rect 3690 1944 3702 1946
rect 3690 1936 3692 1944
rect 3700 1936 3702 1944
rect 3690 1764 3702 1936
rect 3786 1844 3798 1846
rect 3786 1836 3788 1844
rect 3796 1836 3798 1844
rect 3690 1756 3692 1764
rect 3700 1756 3702 1764
rect 3690 1754 3702 1756
rect 3754 1764 3766 1766
rect 3754 1756 3756 1764
rect 3764 1756 3766 1764
rect 3658 1736 3660 1744
rect 3668 1736 3670 1744
rect 3658 1734 3670 1736
rect 3562 1476 3564 1484
rect 3572 1476 3574 1484
rect 3530 1384 3542 1386
rect 3530 1376 3532 1384
rect 3540 1376 3542 1384
rect 3466 1304 3478 1306
rect 3466 1296 3468 1304
rect 3476 1296 3478 1304
rect 3466 1024 3478 1296
rect 3530 1286 3542 1376
rect 3562 1384 3574 1476
rect 3722 1704 3734 1706
rect 3722 1696 3724 1704
rect 3732 1696 3734 1704
rect 3562 1376 3564 1384
rect 3572 1376 3574 1384
rect 3562 1374 3574 1376
rect 3690 1384 3702 1386
rect 3690 1376 3692 1384
rect 3700 1376 3702 1384
rect 3690 1324 3702 1376
rect 3690 1316 3692 1324
rect 3700 1316 3702 1324
rect 3690 1314 3702 1316
rect 3722 1324 3734 1696
rect 3754 1664 3766 1756
rect 3754 1656 3756 1664
rect 3764 1656 3766 1664
rect 3754 1654 3766 1656
rect 3722 1316 3724 1324
rect 3732 1316 3734 1324
rect 3722 1314 3734 1316
rect 3754 1604 3766 1606
rect 3754 1596 3756 1604
rect 3764 1596 3766 1604
rect 3754 1324 3766 1596
rect 3786 1444 3798 1836
rect 3786 1436 3788 1444
rect 3796 1436 3798 1444
rect 3786 1434 3798 1436
rect 3754 1316 3756 1324
rect 3764 1316 3766 1324
rect 3754 1314 3766 1316
rect 3786 1364 3798 1366
rect 3786 1356 3788 1364
rect 3796 1356 3798 1364
rect 3530 1274 3638 1286
rect 3562 1204 3574 1206
rect 3562 1196 3564 1204
rect 3572 1196 3574 1204
rect 3466 1016 3468 1024
rect 3476 1016 3478 1024
rect 3466 1014 3478 1016
rect 3498 1184 3510 1186
rect 3498 1176 3500 1184
rect 3508 1176 3510 1184
rect 3434 896 3436 904
rect 3444 896 3446 904
rect 3434 894 3446 896
rect 3210 876 3212 884
rect 3220 876 3222 884
rect 3210 874 3222 876
rect 3498 744 3510 1176
rect 3498 736 3500 744
rect 3508 736 3510 744
rect 3498 734 3510 736
rect 3530 1144 3542 1146
rect 3530 1136 3532 1144
rect 3540 1136 3542 1144
rect 3530 704 3542 1136
rect 3530 696 3532 704
rect 3540 696 3542 704
rect 3530 694 3542 696
rect 3112 606 3116 614
rect 3124 606 3132 614
rect 3140 606 3148 614
rect 3156 606 3160 614
rect 2794 324 2838 326
rect 2794 316 2828 324
rect 2836 316 2838 324
rect 2794 314 2838 316
rect 2794 304 2806 314
rect 2794 296 2796 304
rect 2804 296 2806 304
rect 2794 294 2806 296
rect 2698 56 2700 64
rect 2708 56 2710 64
rect 2698 54 2710 56
rect 3112 214 3160 606
rect 3274 624 3286 626
rect 3274 616 3276 624
rect 3284 616 3286 624
rect 3274 504 3286 616
rect 3274 496 3276 504
rect 3284 496 3286 504
rect 3274 494 3286 496
rect 3466 584 3478 586
rect 3466 576 3468 584
rect 3476 576 3478 584
rect 3466 464 3478 576
rect 3466 456 3468 464
rect 3476 456 3478 464
rect 3466 454 3478 456
rect 3112 206 3116 214
rect 3124 206 3132 214
rect 3140 206 3148 214
rect 3156 206 3160 214
rect 2602 16 2604 24
rect 2612 16 2614 24
rect 2602 14 2614 16
rect 1560 6 1564 14
rect 1572 6 1580 14
rect 1588 6 1596 14
rect 1604 6 1608 14
rect 1560 -40 1608 6
rect 3112 -40 3160 206
rect 3562 64 3574 1196
rect 3626 1204 3638 1274
rect 3626 1196 3628 1204
rect 3636 1196 3638 1204
rect 3626 1194 3638 1196
rect 3658 1284 3670 1286
rect 3658 1276 3660 1284
rect 3668 1276 3670 1284
rect 3594 1184 3606 1186
rect 3594 1176 3596 1184
rect 3604 1176 3606 1184
rect 3594 904 3606 1176
rect 3658 964 3670 1276
rect 3658 956 3660 964
rect 3668 956 3670 964
rect 3658 954 3670 956
rect 3786 984 3798 1356
rect 3818 1104 3830 1996
rect 3818 1096 3820 1104
rect 3828 1096 3830 1104
rect 3818 1094 3830 1096
rect 3850 1544 3862 2496
rect 3914 2464 3926 2696
rect 4042 2584 4054 2716
rect 4074 2664 4086 3056
rect 4138 2964 4150 3456
rect 4138 2956 4140 2964
rect 4148 2956 4150 2964
rect 4138 2954 4150 2956
rect 4202 3144 4214 3656
rect 4202 3136 4204 3144
rect 4212 3136 4214 3144
rect 4202 2904 4214 3136
rect 4202 2896 4204 2904
rect 4212 2896 4214 2904
rect 4202 2894 4214 2896
rect 4298 2904 4310 2906
rect 4298 2896 4300 2904
rect 4308 2896 4310 2904
rect 4170 2824 4182 2826
rect 4170 2816 4172 2824
rect 4180 2816 4182 2824
rect 4170 2684 4182 2816
rect 4170 2676 4172 2684
rect 4180 2676 4182 2684
rect 4170 2674 4182 2676
rect 4202 2764 4214 2766
rect 4202 2756 4204 2764
rect 4212 2756 4214 2764
rect 4074 2656 4076 2664
rect 4084 2656 4086 2664
rect 4074 2654 4086 2656
rect 4042 2576 4044 2584
rect 4052 2576 4054 2584
rect 4042 2574 4054 2576
rect 4170 2624 4182 2626
rect 4170 2616 4172 2624
rect 4180 2616 4182 2624
rect 3914 2456 3916 2464
rect 3924 2456 3926 2464
rect 3914 2454 3926 2456
rect 4010 2524 4022 2526
rect 4010 2516 4012 2524
rect 4020 2516 4022 2524
rect 3882 2404 3894 2406
rect 3882 2396 3884 2404
rect 3892 2396 3894 2404
rect 3882 1804 3894 2396
rect 3946 2404 3958 2406
rect 3946 2396 3948 2404
rect 3956 2396 3958 2404
rect 3882 1796 3884 1804
rect 3892 1796 3894 1804
rect 3882 1794 3894 1796
rect 3914 2344 3926 2346
rect 3914 2336 3916 2344
rect 3924 2336 3926 2344
rect 3850 1536 3852 1544
rect 3860 1536 3862 1544
rect 3786 976 3788 984
rect 3796 976 3798 984
rect 3594 896 3596 904
rect 3604 896 3606 904
rect 3594 894 3606 896
rect 3722 944 3734 946
rect 3722 936 3724 944
rect 3732 936 3734 944
rect 3722 884 3734 936
rect 3722 876 3724 884
rect 3732 876 3734 884
rect 3722 874 3734 876
rect 3722 724 3734 726
rect 3722 716 3724 724
rect 3732 716 3734 724
rect 3722 686 3734 716
rect 3786 724 3798 976
rect 3786 716 3788 724
rect 3796 716 3798 724
rect 3786 714 3798 716
rect 3818 724 3830 726
rect 3818 716 3820 724
rect 3828 716 3830 724
rect 3818 686 3830 716
rect 3722 674 3830 686
rect 3562 56 3564 64
rect 3572 56 3574 64
rect 3562 54 3574 56
rect 3850 44 3862 1536
rect 3914 1704 3926 2336
rect 3946 2084 3958 2396
rect 3946 2076 3948 2084
rect 3956 2076 3958 2084
rect 3946 2074 3958 2076
rect 4010 2024 4022 2516
rect 4042 2464 4054 2466
rect 4042 2456 4044 2464
rect 4052 2456 4054 2464
rect 4042 2064 4054 2456
rect 4042 2056 4044 2064
rect 4052 2056 4054 2064
rect 4042 2054 4054 2056
rect 4074 2464 4086 2466
rect 4074 2456 4076 2464
rect 4084 2456 4086 2464
rect 4010 2016 4012 2024
rect 4020 2016 4022 2024
rect 4010 2014 4022 2016
rect 3914 1696 3916 1704
rect 3924 1696 3926 1704
rect 3882 1524 3894 1526
rect 3882 1516 3884 1524
rect 3892 1516 3894 1524
rect 3882 1084 3894 1516
rect 3914 1104 3926 1696
rect 3946 1944 3958 1946
rect 3946 1936 3948 1944
rect 3956 1936 3958 1944
rect 3946 1424 3958 1936
rect 4010 1824 4022 1826
rect 4010 1816 4012 1824
rect 4020 1816 4022 1824
rect 3946 1416 3948 1424
rect 3956 1416 3958 1424
rect 3946 1414 3958 1416
rect 3978 1564 3990 1566
rect 3978 1556 3980 1564
rect 3988 1556 3990 1564
rect 3914 1096 3916 1104
rect 3924 1096 3926 1104
rect 3914 1094 3926 1096
rect 3946 1144 3958 1146
rect 3946 1136 3948 1144
rect 3956 1136 3958 1144
rect 3882 1076 3884 1084
rect 3892 1076 3894 1084
rect 3882 1074 3894 1076
rect 3946 1064 3958 1136
rect 3946 1056 3948 1064
rect 3956 1056 3958 1064
rect 3946 1054 3958 1056
rect 3978 1104 3990 1556
rect 3978 1096 3980 1104
rect 3988 1096 3990 1104
rect 3882 984 3894 986
rect 3882 976 3884 984
rect 3892 976 3894 984
rect 3882 404 3894 976
rect 3978 944 3990 1096
rect 4010 984 4022 1816
rect 4042 1644 4054 1646
rect 4042 1636 4044 1644
rect 4052 1636 4054 1644
rect 4042 1344 4054 1636
rect 4042 1336 4044 1344
rect 4052 1336 4054 1344
rect 4042 1334 4054 1336
rect 4010 976 4012 984
rect 4020 976 4022 984
rect 4010 974 4022 976
rect 4042 984 4054 986
rect 4042 976 4044 984
rect 4052 976 4054 984
rect 3978 936 3980 944
rect 3988 936 3990 944
rect 3978 934 3990 936
rect 3882 396 3884 404
rect 3892 396 3894 404
rect 3882 394 3894 396
rect 3914 784 3926 786
rect 3914 776 3916 784
rect 3924 776 3926 784
rect 3914 384 3926 776
rect 3978 744 3990 746
rect 3978 736 3980 744
rect 3988 736 3990 744
rect 3978 564 3990 736
rect 4042 684 4054 976
rect 4042 676 4044 684
rect 4052 676 4054 684
rect 4042 674 4054 676
rect 3978 556 3980 564
rect 3988 556 3990 564
rect 3978 554 3990 556
rect 3914 376 3916 384
rect 3924 376 3926 384
rect 3914 374 3926 376
rect 3978 324 3990 326
rect 3978 316 3980 324
rect 3988 316 3990 324
rect 3978 286 3990 316
rect 3978 284 4022 286
rect 3978 276 4012 284
rect 4020 276 4022 284
rect 3978 274 4022 276
rect 4074 244 4086 2456
rect 4170 2444 4182 2616
rect 4202 2544 4214 2756
rect 4298 2644 4310 2896
rect 4298 2636 4300 2644
rect 4308 2636 4310 2644
rect 4298 2634 4310 2636
rect 4330 2904 4342 2906
rect 4330 2896 4332 2904
rect 4340 2896 4342 2904
rect 4202 2536 4204 2544
rect 4212 2536 4214 2544
rect 4202 2534 4214 2536
rect 4330 2544 4342 2896
rect 4330 2536 4332 2544
rect 4340 2536 4342 2544
rect 4330 2534 4342 2536
rect 4170 2436 4172 2444
rect 4180 2436 4182 2444
rect 4170 2434 4182 2436
rect 4170 2364 4182 2366
rect 4170 2356 4172 2364
rect 4180 2356 4182 2364
rect 4106 2084 4118 2086
rect 4106 2076 4108 2084
rect 4116 2076 4118 2084
rect 4106 1884 4118 2076
rect 4106 1876 4108 1884
rect 4116 1876 4118 1884
rect 4106 1874 4118 1876
rect 4138 2064 4150 2066
rect 4138 2056 4140 2064
rect 4148 2056 4150 2064
rect 4106 1704 4118 1706
rect 4106 1696 4108 1704
rect 4116 1696 4118 1704
rect 4106 1604 4118 1696
rect 4138 1704 4150 2056
rect 4170 1804 4182 2356
rect 4170 1796 4172 1804
rect 4180 1796 4182 1804
rect 4170 1794 4182 1796
rect 4234 1924 4246 1926
rect 4234 1916 4236 1924
rect 4244 1916 4246 1924
rect 4138 1696 4140 1704
rect 4148 1696 4150 1704
rect 4138 1694 4150 1696
rect 4234 1704 4246 1916
rect 4234 1696 4236 1704
rect 4244 1696 4246 1704
rect 4234 1694 4246 1696
rect 4106 1596 4108 1604
rect 4116 1596 4118 1604
rect 4106 1594 4118 1596
rect 4138 1604 4150 1606
rect 4138 1596 4140 1604
rect 4148 1596 4150 1604
rect 4138 1324 4150 1596
rect 4138 1316 4140 1324
rect 4148 1316 4150 1324
rect 4138 1314 4150 1316
rect 4202 1484 4214 1486
rect 4202 1476 4204 1484
rect 4212 1476 4214 1484
rect 4170 1284 4182 1286
rect 4170 1276 4172 1284
rect 4180 1276 4182 1284
rect 4170 964 4182 1276
rect 4170 956 4172 964
rect 4180 956 4182 964
rect 4170 924 4182 956
rect 4170 916 4172 924
rect 4180 916 4182 924
rect 4170 914 4182 916
rect 4074 236 4076 244
rect 4084 236 4086 244
rect 4074 234 4086 236
rect 4170 804 4182 806
rect 4170 796 4172 804
rect 4180 796 4182 804
rect 3850 36 3852 44
rect 3860 36 3862 44
rect 3850 34 3862 36
rect 4170 44 4182 796
rect 4202 804 4214 1476
rect 4362 1264 4374 5156
rect 4586 5084 4598 5336
rect 4586 5076 4588 5084
rect 4596 5076 4598 5084
rect 4586 5074 4598 5076
rect 4632 5214 4680 5606
rect 5226 5644 5238 5646
rect 5226 5636 5228 5644
rect 5236 5636 5238 5644
rect 5194 5544 5206 5546
rect 5194 5536 5196 5544
rect 5204 5536 5206 5544
rect 4632 5206 4636 5214
rect 4644 5206 4652 5214
rect 4660 5206 4668 5214
rect 4676 5206 4680 5214
rect 4458 4944 4470 4946
rect 4458 4936 4460 4944
rect 4468 4936 4470 4944
rect 4394 4744 4406 4746
rect 4394 4736 4396 4744
rect 4404 4736 4406 4744
rect 4394 4604 4406 4736
rect 4394 4596 4396 4604
rect 4404 4596 4406 4604
rect 4394 4594 4406 4596
rect 4458 4444 4470 4936
rect 4632 4814 4680 5206
rect 5130 5264 5142 5266
rect 5130 5256 5132 5264
rect 5140 5256 5142 5264
rect 4632 4806 4636 4814
rect 4644 4806 4652 4814
rect 4660 4806 4668 4814
rect 4676 4806 4680 4814
rect 4586 4504 4598 4506
rect 4586 4496 4588 4504
rect 4596 4496 4598 4504
rect 4458 4436 4460 4444
rect 4468 4436 4470 4444
rect 4458 4434 4470 4436
rect 4490 4464 4502 4466
rect 4490 4456 4492 4464
rect 4500 4456 4502 4464
rect 4458 4284 4470 4286
rect 4458 4276 4460 4284
rect 4468 4276 4470 4284
rect 4458 4084 4470 4276
rect 4490 4104 4502 4456
rect 4586 4244 4598 4496
rect 4586 4236 4588 4244
rect 4596 4236 4598 4244
rect 4586 4234 4598 4236
rect 4632 4414 4680 4806
rect 4906 4944 4918 4946
rect 4906 4936 4908 4944
rect 4916 4936 4918 4944
rect 4906 4904 4918 4936
rect 4906 4896 4908 4904
rect 4916 4896 4918 4904
rect 4906 4504 4918 4896
rect 5130 4884 5142 5256
rect 5194 5104 5206 5536
rect 5194 5096 5196 5104
rect 5204 5096 5206 5104
rect 5194 5094 5206 5096
rect 5130 4876 5132 4884
rect 5140 4876 5142 4884
rect 5130 4874 5142 4876
rect 4906 4496 4908 4504
rect 4916 4496 4918 4504
rect 4906 4494 4918 4496
rect 5002 4764 5014 4766
rect 5002 4756 5004 4764
rect 5012 4756 5014 4764
rect 4632 4406 4636 4414
rect 4644 4406 4652 4414
rect 4660 4406 4668 4414
rect 4676 4406 4680 4414
rect 4490 4096 4492 4104
rect 4500 4096 4502 4104
rect 4490 4094 4502 4096
rect 4458 4076 4460 4084
rect 4468 4076 4470 4084
rect 4458 4074 4470 4076
rect 4632 4014 4680 4406
rect 4746 4204 4758 4206
rect 4746 4196 4748 4204
rect 4756 4196 4758 4204
rect 4746 4064 4758 4196
rect 4746 4056 4748 4064
rect 4756 4056 4758 4064
rect 4746 4054 4758 4056
rect 4874 4124 4886 4126
rect 4874 4116 4876 4124
rect 4884 4116 4886 4124
rect 4874 4044 4886 4116
rect 4874 4036 4876 4044
rect 4884 4036 4886 4044
rect 4874 4034 4886 4036
rect 4632 4006 4636 4014
rect 4644 4006 4652 4014
rect 4660 4006 4668 4014
rect 4676 4006 4680 4014
rect 4586 3924 4598 3926
rect 4586 3916 4588 3924
rect 4596 3916 4598 3924
rect 4458 3644 4470 3646
rect 4458 3636 4460 3644
rect 4468 3636 4470 3644
rect 4458 3084 4470 3636
rect 4458 3076 4460 3084
rect 4468 3076 4470 3084
rect 4458 3074 4470 3076
rect 4490 3344 4502 3346
rect 4490 3336 4492 3344
rect 4500 3336 4502 3344
rect 4490 3084 4502 3336
rect 4490 3076 4492 3084
rect 4500 3076 4502 3084
rect 4490 2984 4502 3076
rect 4586 3064 4598 3916
rect 4586 3056 4588 3064
rect 4596 3056 4598 3064
rect 4586 3054 4598 3056
rect 4632 3614 4680 4006
rect 4632 3606 4636 3614
rect 4644 3606 4652 3614
rect 4660 3606 4668 3614
rect 4676 3606 4680 3614
rect 4632 3214 4680 3606
rect 4746 4004 4758 4006
rect 4746 3996 4748 4004
rect 4756 3996 4758 4004
rect 4746 3524 4758 3996
rect 4746 3516 4748 3524
rect 4756 3516 4758 3524
rect 4746 3514 4758 3516
rect 4632 3206 4636 3214
rect 4644 3206 4652 3214
rect 4660 3206 4668 3214
rect 4676 3206 4680 3214
rect 4490 2976 4492 2984
rect 4500 2976 4502 2984
rect 4490 2726 4502 2976
rect 4554 2884 4566 2886
rect 4554 2876 4556 2884
rect 4564 2876 4566 2884
rect 4490 2714 4534 2726
rect 4490 2384 4502 2386
rect 4490 2376 4492 2384
rect 4500 2376 4502 2384
rect 4394 2324 4406 2326
rect 4394 2316 4396 2324
rect 4404 2316 4406 2324
rect 4394 2044 4406 2316
rect 4490 2304 4502 2376
rect 4490 2296 4492 2304
rect 4500 2296 4502 2304
rect 4490 2294 4502 2296
rect 4394 2036 4396 2044
rect 4404 2036 4406 2044
rect 4394 2034 4406 2036
rect 4426 2204 4438 2206
rect 4426 2196 4428 2204
rect 4436 2196 4438 2204
rect 4426 2044 4438 2196
rect 4426 2036 4428 2044
rect 4436 2036 4438 2044
rect 4426 2034 4438 2036
rect 4522 1864 4534 2714
rect 4554 2444 4566 2876
rect 4632 2814 4680 3206
rect 4632 2806 4636 2814
rect 4644 2806 4652 2814
rect 4660 2806 4668 2814
rect 4676 2806 4680 2814
rect 4554 2436 4556 2444
rect 4564 2436 4566 2444
rect 4554 2434 4566 2436
rect 4586 2704 4598 2706
rect 4586 2696 4588 2704
rect 4596 2696 4598 2704
rect 4586 2524 4598 2696
rect 4586 2516 4588 2524
rect 4596 2516 4598 2524
rect 4586 2304 4598 2516
rect 4586 2296 4588 2304
rect 4596 2296 4598 2304
rect 4586 2294 4598 2296
rect 4632 2414 4680 2806
rect 4842 3324 4854 3326
rect 4842 3316 4844 3324
rect 4852 3316 4854 3324
rect 4632 2406 4636 2414
rect 4644 2406 4652 2414
rect 4660 2406 4668 2414
rect 4676 2406 4680 2414
rect 4554 2284 4566 2286
rect 4554 2276 4556 2284
rect 4564 2276 4566 2284
rect 4554 2124 4566 2276
rect 4554 2116 4556 2124
rect 4564 2116 4566 2124
rect 4554 2114 4566 2116
rect 4522 1856 4524 1864
rect 4532 1856 4534 1864
rect 4522 1854 4534 1856
rect 4632 2014 4680 2406
rect 4714 2764 4726 2766
rect 4714 2756 4716 2764
rect 4724 2756 4726 2764
rect 4714 2064 4726 2756
rect 4778 2724 4790 2726
rect 4778 2716 4780 2724
rect 4788 2716 4790 2724
rect 4778 2444 4790 2716
rect 4778 2436 4780 2444
rect 4788 2436 4790 2444
rect 4778 2434 4790 2436
rect 4810 2704 4822 2706
rect 4810 2696 4812 2704
rect 4820 2696 4822 2704
rect 4810 2284 4822 2696
rect 4810 2276 4812 2284
rect 4820 2276 4822 2284
rect 4810 2274 4822 2276
rect 4842 2104 4854 3316
rect 4906 3304 4918 3306
rect 4906 3296 4908 3304
rect 4916 3296 4918 3304
rect 4842 2096 4844 2104
rect 4852 2096 4854 2104
rect 4842 2094 4854 2096
rect 4874 2444 4886 2446
rect 4874 2436 4876 2444
rect 4884 2436 4886 2444
rect 4714 2056 4716 2064
rect 4724 2056 4726 2064
rect 4714 2054 4726 2056
rect 4746 2064 4758 2066
rect 4746 2056 4748 2064
rect 4756 2056 4758 2064
rect 4746 2024 4758 2056
rect 4746 2016 4748 2024
rect 4756 2016 4758 2024
rect 4746 2014 4758 2016
rect 4632 2006 4636 2014
rect 4644 2006 4652 2014
rect 4660 2006 4668 2014
rect 4676 2006 4680 2014
rect 4632 1614 4680 2006
rect 4810 2004 4822 2006
rect 4810 1996 4812 2004
rect 4820 1996 4822 2004
rect 4810 1904 4822 1996
rect 4810 1896 4812 1904
rect 4820 1896 4822 1904
rect 4810 1894 4822 1896
rect 4842 2004 4854 2006
rect 4842 1996 4844 2004
rect 4852 1996 4854 2004
rect 4714 1864 4726 1866
rect 4714 1856 4716 1864
rect 4724 1856 4726 1864
rect 4714 1804 4726 1856
rect 4714 1796 4716 1804
rect 4724 1796 4726 1804
rect 4714 1794 4726 1796
rect 4632 1606 4636 1614
rect 4644 1606 4652 1614
rect 4660 1606 4668 1614
rect 4676 1606 4680 1614
rect 4458 1484 4470 1486
rect 4458 1476 4460 1484
rect 4468 1476 4470 1484
rect 4426 1344 4438 1346
rect 4426 1336 4428 1344
rect 4436 1336 4438 1344
rect 4362 1256 4364 1264
rect 4372 1256 4374 1264
rect 4362 1254 4374 1256
rect 4394 1264 4406 1266
rect 4394 1256 4396 1264
rect 4404 1256 4406 1264
rect 4202 796 4204 804
rect 4212 796 4214 804
rect 4202 794 4214 796
rect 4330 1224 4342 1226
rect 4330 1216 4332 1224
rect 4340 1216 4342 1224
rect 4330 784 4342 1216
rect 4394 944 4406 1256
rect 4426 1204 4438 1336
rect 4426 1196 4428 1204
rect 4436 1196 4438 1204
rect 4426 1194 4438 1196
rect 4394 936 4396 944
rect 4404 936 4406 944
rect 4394 934 4406 936
rect 4458 824 4470 1476
rect 4554 1384 4566 1386
rect 4554 1376 4556 1384
rect 4564 1376 4566 1384
rect 4554 1084 4566 1376
rect 4554 1076 4556 1084
rect 4564 1076 4566 1084
rect 4554 1074 4566 1076
rect 4632 1214 4680 1606
rect 4778 1764 4790 1766
rect 4778 1756 4780 1764
rect 4788 1756 4790 1764
rect 4778 1504 4790 1756
rect 4778 1496 4780 1504
rect 4788 1496 4790 1504
rect 4778 1494 4790 1496
rect 4810 1564 4822 1566
rect 4810 1556 4812 1564
rect 4820 1556 4822 1564
rect 4632 1206 4636 1214
rect 4644 1206 4652 1214
rect 4660 1206 4668 1214
rect 4676 1206 4680 1214
rect 4458 816 4460 824
rect 4468 816 4470 824
rect 4458 814 4470 816
rect 4554 1004 4566 1006
rect 4554 996 4556 1004
rect 4564 996 4566 1004
rect 4330 776 4332 784
rect 4340 776 4342 784
rect 4330 774 4342 776
rect 4522 624 4534 626
rect 4522 616 4524 624
rect 4532 616 4534 624
rect 4522 524 4534 616
rect 4522 516 4524 524
rect 4532 516 4534 524
rect 4522 514 4534 516
rect 4554 324 4566 996
rect 4554 316 4556 324
rect 4564 316 4566 324
rect 4554 314 4566 316
rect 4632 814 4680 1206
rect 4632 806 4636 814
rect 4644 806 4652 814
rect 4660 806 4668 814
rect 4676 806 4680 814
rect 4632 414 4680 806
rect 4632 406 4636 414
rect 4644 406 4652 414
rect 4660 406 4668 414
rect 4676 406 4680 414
rect 4170 36 4172 44
rect 4180 36 4182 44
rect 4170 34 4182 36
rect 4632 14 4680 406
rect 4746 684 4758 686
rect 4746 676 4748 684
rect 4756 676 4758 684
rect 4746 404 4758 676
rect 4746 396 4748 404
rect 4756 396 4758 404
rect 4746 394 4758 396
rect 4810 24 4822 1556
rect 4842 1264 4854 1996
rect 4874 1704 4886 2436
rect 4906 2344 4918 3296
rect 5002 3024 5014 4756
rect 5130 4544 5142 4546
rect 5130 4536 5132 4544
rect 5140 4536 5142 4544
rect 5130 4264 5142 4536
rect 5226 4544 5238 5636
rect 5546 5584 5558 5586
rect 5546 5576 5548 5584
rect 5556 5576 5558 5584
rect 5450 5524 5462 5526
rect 5450 5516 5452 5524
rect 5460 5516 5462 5524
rect 5450 5486 5462 5516
rect 5386 5474 5462 5486
rect 5386 5464 5398 5474
rect 5386 5456 5388 5464
rect 5396 5456 5398 5464
rect 5386 5454 5398 5456
rect 5226 4536 5228 4544
rect 5236 4536 5238 4544
rect 5226 4534 5238 4536
rect 5258 4924 5270 4926
rect 5258 4916 5260 4924
rect 5268 4916 5270 4924
rect 5258 4524 5270 4916
rect 5258 4516 5260 4524
rect 5268 4516 5270 4524
rect 5130 4256 5132 4264
rect 5140 4256 5142 4264
rect 5130 4254 5142 4256
rect 5162 4344 5174 4346
rect 5162 4336 5164 4344
rect 5172 4336 5174 4344
rect 5162 4304 5174 4336
rect 5162 4296 5164 4304
rect 5172 4296 5174 4304
rect 5162 4124 5174 4296
rect 5162 4116 5164 4124
rect 5172 4116 5174 4124
rect 5162 4114 5174 4116
rect 5162 4064 5174 4066
rect 5162 4056 5164 4064
rect 5172 4056 5174 4064
rect 5130 3804 5142 3806
rect 5130 3796 5132 3804
rect 5140 3796 5142 3804
rect 5066 3424 5078 3426
rect 5066 3416 5068 3424
rect 5076 3416 5078 3424
rect 5066 3344 5078 3416
rect 5066 3336 5068 3344
rect 5076 3336 5078 3344
rect 5066 3334 5078 3336
rect 5002 3016 5004 3024
rect 5012 3016 5014 3024
rect 5002 3014 5014 3016
rect 5098 2964 5110 2966
rect 5098 2956 5100 2964
rect 5108 2956 5110 2964
rect 5034 2924 5046 2926
rect 5034 2916 5036 2924
rect 5044 2916 5046 2924
rect 4970 2884 4982 2886
rect 4970 2876 4972 2884
rect 4980 2876 4982 2884
rect 4906 2336 4908 2344
rect 4916 2336 4918 2344
rect 4906 2334 4918 2336
rect 4938 2644 4950 2646
rect 4938 2636 4940 2644
rect 4948 2636 4950 2644
rect 4938 2284 4950 2636
rect 4970 2484 4982 2876
rect 5034 2544 5046 2916
rect 5034 2536 5036 2544
rect 5044 2536 5046 2544
rect 5034 2534 5046 2536
rect 5066 2764 5078 2766
rect 5066 2756 5068 2764
rect 5076 2756 5078 2764
rect 4970 2476 4972 2484
rect 4980 2476 4982 2484
rect 4970 2474 4982 2476
rect 4938 2276 4940 2284
rect 4948 2276 4950 2284
rect 4938 2274 4950 2276
rect 4970 2384 4982 2386
rect 4970 2376 4972 2384
rect 4980 2376 4982 2384
rect 4970 2064 4982 2376
rect 4970 2056 4972 2064
rect 4980 2056 4982 2064
rect 4970 2054 4982 2056
rect 5066 1984 5078 2756
rect 5098 2764 5110 2956
rect 5098 2756 5100 2764
rect 5108 2756 5110 2764
rect 5098 2754 5110 2756
rect 5098 2724 5110 2726
rect 5098 2716 5100 2724
rect 5108 2716 5110 2724
rect 5098 2384 5110 2716
rect 5130 2724 5142 3796
rect 5162 3184 5174 4056
rect 5258 3904 5270 4516
rect 5290 4804 5302 4806
rect 5290 4796 5292 4804
rect 5300 4796 5302 4804
rect 5290 4524 5302 4796
rect 5290 4516 5292 4524
rect 5300 4516 5302 4524
rect 5290 4514 5302 4516
rect 5386 4664 5398 4666
rect 5386 4656 5388 4664
rect 5396 4656 5398 4664
rect 5386 4504 5398 4656
rect 5386 4496 5388 4504
rect 5396 4496 5398 4504
rect 5354 4324 5366 4326
rect 5354 4316 5356 4324
rect 5364 4316 5366 4324
rect 5258 3896 5260 3904
rect 5268 3896 5270 3904
rect 5258 3894 5270 3896
rect 5290 4264 5302 4266
rect 5290 4256 5292 4264
rect 5300 4256 5302 4264
rect 5290 3884 5302 4256
rect 5354 4164 5366 4316
rect 5386 4204 5398 4496
rect 5514 4644 5526 4646
rect 5514 4636 5516 4644
rect 5524 4636 5526 4644
rect 5386 4196 5388 4204
rect 5396 4196 5398 4204
rect 5386 4194 5398 4196
rect 5450 4284 5462 4286
rect 5450 4276 5452 4284
rect 5460 4276 5462 4284
rect 5450 4204 5462 4276
rect 5450 4196 5452 4204
rect 5460 4196 5462 4204
rect 5450 4194 5462 4196
rect 5354 4156 5356 4164
rect 5364 4156 5366 4164
rect 5354 4154 5366 4156
rect 5450 4124 5462 4126
rect 5450 4116 5452 4124
rect 5460 4116 5462 4124
rect 5418 4084 5430 4086
rect 5418 4076 5420 4084
rect 5428 4076 5430 4084
rect 5386 4044 5398 4046
rect 5386 4036 5388 4044
rect 5396 4036 5398 4044
rect 5354 3964 5366 3966
rect 5354 3956 5356 3964
rect 5364 3956 5366 3964
rect 5290 3876 5292 3884
rect 5300 3876 5302 3884
rect 5290 3874 5302 3876
rect 5322 3904 5334 3906
rect 5322 3896 5324 3904
rect 5332 3896 5334 3904
rect 5322 3846 5334 3896
rect 5274 3844 5334 3846
rect 5274 3836 5276 3844
rect 5284 3836 5334 3844
rect 5274 3834 5334 3836
rect 5290 3784 5302 3786
rect 5290 3776 5292 3784
rect 5300 3776 5302 3784
rect 5162 3176 5164 3184
rect 5172 3176 5174 3184
rect 5162 3174 5174 3176
rect 5226 3724 5238 3726
rect 5226 3716 5228 3724
rect 5236 3716 5238 3724
rect 5130 2716 5132 2724
rect 5140 2716 5142 2724
rect 5130 2714 5142 2716
rect 5162 3024 5174 3026
rect 5162 3016 5164 3024
rect 5172 3016 5174 3024
rect 5130 2624 5142 2626
rect 5130 2616 5132 2624
rect 5140 2616 5142 2624
rect 5130 2504 5142 2616
rect 5130 2496 5132 2504
rect 5140 2496 5142 2504
rect 5130 2494 5142 2496
rect 5098 2376 5100 2384
rect 5108 2376 5110 2384
rect 5098 2374 5110 2376
rect 5098 2344 5110 2346
rect 5098 2336 5100 2344
rect 5108 2336 5110 2344
rect 5098 2144 5110 2336
rect 5098 2136 5100 2144
rect 5108 2136 5110 2144
rect 5098 2134 5110 2136
rect 5130 2284 5142 2286
rect 5130 2276 5132 2284
rect 5140 2276 5142 2284
rect 5130 2044 5142 2276
rect 5162 2064 5174 3016
rect 5226 2544 5238 3716
rect 5258 3444 5270 3446
rect 5258 3436 5260 3444
rect 5268 3436 5270 3444
rect 5258 2964 5270 3436
rect 5290 3444 5302 3776
rect 5290 3436 5292 3444
rect 5300 3436 5302 3444
rect 5290 3434 5302 3436
rect 5258 2956 5260 2964
rect 5268 2956 5270 2964
rect 5258 2954 5270 2956
rect 5290 3024 5302 3026
rect 5290 3016 5292 3024
rect 5300 3016 5302 3024
rect 5226 2536 5228 2544
rect 5236 2536 5238 2544
rect 5226 2534 5238 2536
rect 5258 2924 5270 2926
rect 5258 2916 5260 2924
rect 5268 2916 5270 2924
rect 5258 2544 5270 2916
rect 5258 2536 5260 2544
rect 5268 2536 5270 2544
rect 5258 2534 5270 2536
rect 5162 2056 5164 2064
rect 5172 2056 5174 2064
rect 5162 2054 5174 2056
rect 5258 2384 5270 2386
rect 5258 2376 5260 2384
rect 5268 2376 5270 2384
rect 5130 2036 5132 2044
rect 5140 2036 5142 2044
rect 5130 2034 5142 2036
rect 5066 1976 5068 1984
rect 5076 1976 5078 1984
rect 5066 1974 5078 1976
rect 5194 1804 5206 1806
rect 5194 1796 5196 1804
rect 5204 1796 5206 1804
rect 4874 1696 4876 1704
rect 4884 1696 4886 1704
rect 4874 1694 4886 1696
rect 5034 1784 5046 1786
rect 5034 1776 5036 1784
rect 5044 1776 5046 1784
rect 5034 1364 5046 1776
rect 5034 1356 5036 1364
rect 5044 1356 5046 1364
rect 5034 1354 5046 1356
rect 4842 1256 4844 1264
rect 4852 1256 4854 1264
rect 4842 1254 4854 1256
rect 4970 1344 4982 1346
rect 4970 1336 4972 1344
rect 4980 1336 4982 1344
rect 4970 944 4982 1336
rect 5194 1344 5206 1796
rect 5258 1604 5270 2376
rect 5290 2324 5302 3016
rect 5290 2316 5292 2324
rect 5300 2316 5302 2324
rect 5290 2314 5302 2316
rect 5322 2964 5334 2966
rect 5322 2956 5324 2964
rect 5332 2956 5334 2964
rect 5258 1596 5260 1604
rect 5268 1596 5270 1604
rect 5258 1594 5270 1596
rect 5194 1336 5196 1344
rect 5204 1336 5206 1344
rect 5194 1334 5206 1336
rect 4970 936 4972 944
rect 4980 936 4982 944
rect 4970 934 4982 936
rect 5034 1104 5046 1106
rect 5034 1096 5036 1104
rect 5044 1096 5046 1104
rect 5034 724 5046 1096
rect 5258 1084 5270 1086
rect 5258 1076 5260 1084
rect 5268 1076 5270 1084
rect 5130 1004 5142 1006
rect 5130 996 5132 1004
rect 5140 996 5142 1004
rect 5130 944 5142 996
rect 5130 936 5132 944
rect 5140 936 5142 944
rect 5130 934 5142 936
rect 5034 716 5036 724
rect 5044 716 5046 724
rect 5034 714 5046 716
rect 5258 664 5270 1076
rect 5322 824 5334 2956
rect 5354 2964 5366 3956
rect 5386 3024 5398 4036
rect 5418 3144 5430 4076
rect 5418 3136 5420 3144
rect 5428 3136 5430 3144
rect 5418 3134 5430 3136
rect 5450 4024 5462 4116
rect 5450 4016 5452 4024
rect 5460 4016 5462 4024
rect 5450 3084 5462 4016
rect 5482 4084 5494 4086
rect 5482 4076 5484 4084
rect 5492 4076 5494 4084
rect 5482 3244 5494 4076
rect 5514 4044 5526 4636
rect 5514 4036 5516 4044
rect 5524 4036 5526 4044
rect 5514 4034 5526 4036
rect 5514 3724 5526 3726
rect 5514 3716 5516 3724
rect 5524 3716 5526 3724
rect 5514 3324 5526 3716
rect 5546 3504 5558 5576
rect 5642 5404 5654 5406
rect 5642 5396 5644 5404
rect 5652 5396 5654 5404
rect 5578 5224 5590 5226
rect 5578 5216 5580 5224
rect 5588 5216 5590 5224
rect 5578 4344 5590 5216
rect 5642 4524 5654 5396
rect 5898 5404 5910 5736
rect 5898 5396 5900 5404
rect 5908 5396 5910 5404
rect 5898 5394 5910 5396
rect 6026 5684 6038 5686
rect 6026 5676 6028 5684
rect 6036 5676 6038 5684
rect 5834 5344 5846 5346
rect 5834 5336 5836 5344
rect 5844 5336 5846 5344
rect 5642 4516 5644 4524
rect 5652 4516 5654 4524
rect 5642 4514 5654 4516
rect 5738 5144 5750 5146
rect 5738 5136 5740 5144
rect 5748 5136 5750 5144
rect 5578 4336 5580 4344
rect 5588 4336 5590 4344
rect 5578 4334 5590 4336
rect 5706 4424 5718 4426
rect 5706 4416 5708 4424
rect 5716 4416 5718 4424
rect 5642 4304 5654 4306
rect 5642 4296 5644 4304
rect 5652 4296 5654 4304
rect 5642 4184 5654 4296
rect 5706 4244 5718 4416
rect 5738 4384 5750 5136
rect 5738 4376 5740 4384
rect 5748 4376 5750 4384
rect 5738 4374 5750 4376
rect 5770 5044 5782 5046
rect 5770 5036 5772 5044
rect 5780 5036 5782 5044
rect 5706 4236 5708 4244
rect 5716 4236 5718 4244
rect 5706 4234 5718 4236
rect 5738 4324 5750 4326
rect 5738 4316 5740 4324
rect 5748 4316 5750 4324
rect 5738 4244 5750 4316
rect 5738 4236 5740 4244
rect 5748 4236 5750 4244
rect 5642 4176 5644 4184
rect 5652 4176 5654 4184
rect 5642 4174 5654 4176
rect 5674 4144 5686 4146
rect 5674 4136 5676 4144
rect 5684 4136 5686 4144
rect 5642 4104 5654 4106
rect 5642 4096 5644 4104
rect 5652 4096 5654 4104
rect 5610 3864 5622 3866
rect 5610 3856 5612 3864
rect 5620 3856 5622 3864
rect 5610 3744 5622 3856
rect 5642 3784 5654 4096
rect 5674 4084 5686 4136
rect 5674 4076 5676 4084
rect 5684 4076 5686 4084
rect 5674 4074 5686 4076
rect 5642 3776 5644 3784
rect 5652 3776 5654 3784
rect 5642 3774 5654 3776
rect 5706 3924 5718 3926
rect 5706 3916 5708 3924
rect 5716 3916 5718 3924
rect 5610 3736 5612 3744
rect 5620 3736 5622 3744
rect 5610 3734 5622 3736
rect 5546 3496 5548 3504
rect 5556 3496 5558 3504
rect 5546 3494 5558 3496
rect 5642 3704 5654 3706
rect 5642 3696 5644 3704
rect 5652 3696 5654 3704
rect 5514 3316 5516 3324
rect 5524 3316 5526 3324
rect 5514 3314 5526 3316
rect 5578 3404 5590 3406
rect 5578 3396 5580 3404
rect 5588 3396 5590 3404
rect 5482 3236 5484 3244
rect 5492 3236 5494 3244
rect 5482 3234 5494 3236
rect 5450 3076 5452 3084
rect 5460 3076 5462 3084
rect 5450 3074 5462 3076
rect 5386 3016 5388 3024
rect 5396 3016 5398 3024
rect 5386 3014 5398 3016
rect 5354 2956 5356 2964
rect 5364 2956 5366 2964
rect 5354 2954 5366 2956
rect 5514 2964 5526 2966
rect 5514 2956 5516 2964
rect 5524 2956 5526 2964
rect 5386 2924 5398 2926
rect 5386 2916 5388 2924
rect 5396 2916 5398 2924
rect 5354 2904 5366 2906
rect 5354 2896 5356 2904
rect 5364 2896 5366 2904
rect 5354 2564 5366 2896
rect 5354 2556 5356 2564
rect 5364 2556 5366 2564
rect 5354 2554 5366 2556
rect 5386 2524 5398 2916
rect 5386 2516 5388 2524
rect 5396 2516 5398 2524
rect 5386 2514 5398 2516
rect 5418 2824 5430 2826
rect 5418 2816 5420 2824
rect 5428 2816 5430 2824
rect 5386 2384 5398 2386
rect 5386 2376 5388 2384
rect 5396 2376 5398 2384
rect 5354 2324 5366 2326
rect 5354 2316 5356 2324
rect 5364 2316 5366 2324
rect 5354 1264 5366 2316
rect 5386 1564 5398 2376
rect 5418 2364 5430 2816
rect 5482 2764 5494 2766
rect 5482 2756 5484 2764
rect 5492 2756 5494 2764
rect 5482 2726 5494 2756
rect 5450 2714 5494 2726
rect 5450 2664 5462 2714
rect 5450 2656 5452 2664
rect 5460 2656 5462 2664
rect 5450 2654 5462 2656
rect 5482 2664 5494 2666
rect 5482 2656 5484 2664
rect 5492 2656 5494 2664
rect 5418 2356 5420 2364
rect 5428 2356 5430 2364
rect 5418 2354 5430 2356
rect 5482 2324 5494 2656
rect 5482 2316 5484 2324
rect 5492 2316 5494 2324
rect 5482 2314 5494 2316
rect 5386 1556 5388 1564
rect 5396 1556 5398 1564
rect 5386 1554 5398 1556
rect 5418 2284 5430 2286
rect 5418 2276 5420 2284
rect 5428 2276 5430 2284
rect 5354 1256 5356 1264
rect 5364 1256 5366 1264
rect 5354 1254 5366 1256
rect 5322 816 5324 824
rect 5332 816 5334 824
rect 5322 814 5334 816
rect 5258 656 5260 664
rect 5268 656 5270 664
rect 5258 654 5270 656
rect 5354 804 5366 806
rect 5354 796 5356 804
rect 5364 796 5366 804
rect 5066 644 5078 646
rect 5066 636 5068 644
rect 5076 636 5078 644
rect 5066 284 5078 636
rect 5066 276 5068 284
rect 5076 276 5078 284
rect 5066 274 5078 276
rect 5354 244 5366 796
rect 5386 584 5398 586
rect 5386 576 5388 584
rect 5396 576 5398 584
rect 5386 324 5398 576
rect 5418 464 5430 2276
rect 5482 2164 5494 2166
rect 5482 2156 5484 2164
rect 5492 2156 5494 2164
rect 5482 844 5494 2156
rect 5514 1944 5526 2956
rect 5578 2924 5590 3396
rect 5578 2916 5580 2924
rect 5588 2916 5590 2924
rect 5578 2914 5590 2916
rect 5642 2904 5654 3696
rect 5642 2896 5644 2904
rect 5652 2896 5654 2904
rect 5642 2894 5654 2896
rect 5674 3384 5686 3386
rect 5674 3376 5676 3384
rect 5684 3376 5686 3384
rect 5514 1936 5516 1944
rect 5524 1936 5526 1944
rect 5514 1934 5526 1936
rect 5546 2864 5558 2866
rect 5546 2856 5548 2864
rect 5556 2856 5558 2864
rect 5546 1684 5558 2856
rect 5642 2864 5654 2866
rect 5642 2856 5644 2864
rect 5652 2856 5654 2864
rect 5610 2644 5622 2646
rect 5610 2636 5612 2644
rect 5620 2636 5622 2644
rect 5578 2624 5590 2626
rect 5578 2616 5580 2624
rect 5588 2616 5590 2624
rect 5578 2384 5590 2616
rect 5578 2376 5580 2384
rect 5588 2376 5590 2384
rect 5578 2374 5590 2376
rect 5610 2284 5622 2636
rect 5610 2276 5612 2284
rect 5620 2276 5622 2284
rect 5610 2274 5622 2276
rect 5642 2244 5654 2856
rect 5674 2544 5686 3376
rect 5706 3324 5718 3916
rect 5706 3316 5708 3324
rect 5716 3316 5718 3324
rect 5706 3314 5718 3316
rect 5706 3284 5718 3286
rect 5706 3276 5708 3284
rect 5716 3276 5718 3284
rect 5706 3104 5718 3276
rect 5738 3284 5750 4236
rect 5738 3276 5740 3284
rect 5748 3276 5750 3284
rect 5738 3274 5750 3276
rect 5706 3096 5708 3104
rect 5716 3096 5718 3104
rect 5706 3094 5718 3096
rect 5738 3124 5750 3126
rect 5738 3116 5740 3124
rect 5748 3116 5750 3124
rect 5674 2536 5676 2544
rect 5684 2536 5686 2544
rect 5674 2534 5686 2536
rect 5706 2964 5718 2966
rect 5706 2956 5708 2964
rect 5716 2956 5718 2964
rect 5642 2236 5644 2244
rect 5652 2236 5654 2244
rect 5642 2234 5654 2236
rect 5706 2184 5718 2956
rect 5738 2864 5750 3116
rect 5770 3064 5782 5036
rect 5802 4344 5814 4346
rect 5802 4336 5804 4344
rect 5812 4336 5814 4344
rect 5802 4144 5814 4336
rect 5802 4136 5804 4144
rect 5812 4136 5814 4144
rect 5802 4134 5814 4136
rect 5770 3056 5772 3064
rect 5780 3056 5782 3064
rect 5770 3054 5782 3056
rect 5802 3744 5814 3746
rect 5802 3736 5804 3744
rect 5812 3736 5814 3744
rect 5738 2856 5740 2864
rect 5748 2856 5750 2864
rect 5738 2854 5750 2856
rect 5770 3024 5782 3026
rect 5770 3016 5772 3024
rect 5780 3016 5782 3024
rect 5738 2744 5750 2746
rect 5738 2736 5740 2744
rect 5748 2736 5750 2744
rect 5738 2644 5750 2736
rect 5738 2636 5740 2644
rect 5748 2636 5750 2644
rect 5738 2634 5750 2636
rect 5738 2344 5750 2346
rect 5738 2336 5740 2344
rect 5748 2336 5750 2344
rect 5738 2204 5750 2336
rect 5738 2196 5740 2204
rect 5748 2196 5750 2204
rect 5738 2194 5750 2196
rect 5706 2176 5708 2184
rect 5716 2176 5718 2184
rect 5706 2174 5718 2176
rect 5610 2164 5622 2166
rect 5610 2156 5612 2164
rect 5620 2156 5622 2164
rect 5610 2024 5622 2156
rect 5610 2016 5612 2024
rect 5620 2016 5622 2024
rect 5610 2014 5622 2016
rect 5706 1944 5718 1946
rect 5706 1936 5708 1944
rect 5716 1936 5718 1944
rect 5706 1926 5718 1936
rect 5642 1924 5718 1926
rect 5642 1916 5644 1924
rect 5652 1916 5718 1924
rect 5642 1914 5718 1916
rect 5546 1676 5548 1684
rect 5556 1676 5558 1684
rect 5482 836 5484 844
rect 5492 836 5494 844
rect 5482 834 5494 836
rect 5514 1044 5526 1046
rect 5514 1036 5516 1044
rect 5524 1036 5526 1044
rect 5514 724 5526 1036
rect 5514 716 5516 724
rect 5524 716 5526 724
rect 5514 714 5526 716
rect 5418 456 5420 464
rect 5428 456 5430 464
rect 5418 454 5430 456
rect 5386 316 5388 324
rect 5396 316 5398 324
rect 5386 314 5398 316
rect 5546 324 5558 1676
rect 5770 1484 5782 3016
rect 5802 2944 5814 3736
rect 5802 2936 5804 2944
rect 5812 2936 5814 2944
rect 5802 2934 5814 2936
rect 5834 3084 5846 5336
rect 5930 5324 5942 5326
rect 5930 5316 5932 5324
rect 5940 5316 5942 5324
rect 5930 4744 5942 5316
rect 5962 5124 5974 5126
rect 5962 5116 5964 5124
rect 5972 5116 5974 5124
rect 5962 4984 5974 5116
rect 5962 4976 5964 4984
rect 5972 4976 5974 4984
rect 5962 4974 5974 4976
rect 6026 4944 6038 5676
rect 6250 5544 6262 5546
rect 6250 5536 6252 5544
rect 6260 5536 6262 5544
rect 6090 5504 6102 5506
rect 6090 5496 6092 5504
rect 6100 5496 6102 5504
rect 6026 4936 6028 4944
rect 6036 4936 6038 4944
rect 6026 4934 6038 4936
rect 6058 5064 6070 5066
rect 6058 5056 6060 5064
rect 6068 5056 6070 5064
rect 5930 4736 5932 4744
rect 5940 4736 5942 4744
rect 5930 4734 5942 4736
rect 5962 4924 5974 4926
rect 5962 4916 5964 4924
rect 5972 4916 5974 4924
rect 5834 3076 5836 3084
rect 5844 3076 5846 3084
rect 5802 2864 5814 2866
rect 5802 2856 5804 2864
rect 5812 2856 5814 2864
rect 5802 2504 5814 2856
rect 5802 2496 5804 2504
rect 5812 2496 5814 2504
rect 5802 2494 5814 2496
rect 5802 2384 5814 2386
rect 5802 2376 5804 2384
rect 5812 2376 5814 2384
rect 5802 2304 5814 2376
rect 5802 2296 5804 2304
rect 5812 2296 5814 2304
rect 5802 2294 5814 2296
rect 5770 1476 5772 1484
rect 5780 1476 5782 1484
rect 5770 1474 5782 1476
rect 5802 1804 5814 1806
rect 5802 1796 5804 1804
rect 5812 1796 5814 1804
rect 5642 1364 5654 1366
rect 5642 1356 5644 1364
rect 5652 1356 5654 1364
rect 5578 744 5590 746
rect 5578 736 5580 744
rect 5588 736 5590 744
rect 5578 344 5590 736
rect 5578 336 5580 344
rect 5588 336 5590 344
rect 5578 334 5590 336
rect 5546 316 5548 324
rect 5556 316 5558 324
rect 5546 314 5558 316
rect 5354 236 5356 244
rect 5364 236 5366 244
rect 5354 234 5366 236
rect 5418 124 5462 126
rect 5418 116 5420 124
rect 5428 116 5462 124
rect 5418 114 5462 116
rect 5450 104 5462 114
rect 5450 96 5452 104
rect 5460 96 5462 104
rect 5450 94 5462 96
rect 5642 104 5654 1356
rect 5802 124 5814 1796
rect 5834 1744 5846 3076
rect 5834 1736 5836 1744
rect 5844 1736 5846 1744
rect 5834 1734 5846 1736
rect 5866 4704 5878 4706
rect 5866 4696 5868 4704
rect 5876 4696 5878 4704
rect 5834 1704 5846 1706
rect 5834 1696 5836 1704
rect 5844 1696 5846 1704
rect 5834 304 5846 1696
rect 5866 1684 5878 4696
rect 5898 4664 5910 4666
rect 5898 4656 5900 4664
rect 5908 4656 5910 4664
rect 5898 3704 5910 4656
rect 5930 4484 5942 4486
rect 5930 4476 5932 4484
rect 5940 4476 5942 4484
rect 5930 3804 5942 4476
rect 5962 4264 5974 4916
rect 6026 4884 6038 4886
rect 6026 4876 6028 4884
rect 6036 4876 6038 4884
rect 6026 4444 6038 4876
rect 6026 4436 6028 4444
rect 6036 4436 6038 4444
rect 6026 4434 6038 4436
rect 5962 4256 5964 4264
rect 5972 4256 5974 4264
rect 5962 4254 5974 4256
rect 6026 4364 6038 4366
rect 6026 4356 6028 4364
rect 6036 4356 6038 4364
rect 5930 3796 5932 3804
rect 5940 3796 5942 3804
rect 5930 3794 5942 3796
rect 5962 4204 5974 4206
rect 5962 4196 5964 4204
rect 5972 4196 5974 4204
rect 5898 3696 5900 3704
rect 5908 3696 5910 3704
rect 5898 3694 5910 3696
rect 5930 3704 5942 3706
rect 5930 3696 5932 3704
rect 5940 3696 5942 3704
rect 5930 3544 5942 3696
rect 5930 3536 5932 3544
rect 5940 3536 5942 3544
rect 5930 3534 5942 3536
rect 5898 3324 5910 3326
rect 5898 3316 5900 3324
rect 5908 3316 5910 3324
rect 5898 2724 5910 3316
rect 5962 3324 5974 4196
rect 6026 4166 6038 4356
rect 5994 4154 6038 4166
rect 5994 4064 6006 4154
rect 5994 4056 5996 4064
rect 6004 4056 6006 4064
rect 5994 4054 6006 4056
rect 6026 3744 6038 3746
rect 6026 3736 6028 3744
rect 6036 3736 6038 3744
rect 5962 3316 5964 3324
rect 5972 3316 5974 3324
rect 5962 3314 5974 3316
rect 5994 3684 6006 3686
rect 5994 3676 5996 3684
rect 6004 3676 6006 3684
rect 5962 3204 5974 3206
rect 5962 3196 5964 3204
rect 5972 3196 5974 3204
rect 5962 3044 5974 3196
rect 5994 3164 6006 3676
rect 6026 3224 6038 3736
rect 6058 3584 6070 5056
rect 6090 4704 6102 5496
rect 6154 5484 6166 5486
rect 6154 5476 6156 5484
rect 6164 5476 6166 5484
rect 6090 4696 6092 4704
rect 6100 4696 6102 4704
rect 6090 4694 6102 4696
rect 6122 5324 6134 5326
rect 6122 5316 6124 5324
rect 6132 5316 6134 5324
rect 6122 4984 6134 5316
rect 6122 4976 6124 4984
rect 6132 4976 6134 4984
rect 6122 4544 6134 4976
rect 6154 4664 6166 5476
rect 6218 5344 6230 5346
rect 6218 5336 6220 5344
rect 6228 5336 6230 5344
rect 6218 5304 6230 5336
rect 6218 5296 6220 5304
rect 6228 5296 6230 5304
rect 6154 4656 6156 4664
rect 6164 4656 6166 4664
rect 6154 4654 6166 4656
rect 6186 5244 6198 5246
rect 6186 5236 6188 5244
rect 6196 5236 6198 5244
rect 6122 4536 6124 4544
rect 6132 4536 6134 4544
rect 6122 4534 6134 4536
rect 6154 4544 6166 4546
rect 6154 4536 6156 4544
rect 6164 4536 6166 4544
rect 6122 4444 6134 4446
rect 6122 4436 6124 4444
rect 6132 4436 6134 4444
rect 6090 4344 6102 4346
rect 6090 4336 6092 4344
rect 6100 4336 6102 4344
rect 6090 4184 6102 4336
rect 6122 4284 6134 4436
rect 6122 4276 6124 4284
rect 6132 4276 6134 4284
rect 6122 4274 6134 4276
rect 6090 4176 6092 4184
rect 6100 4176 6102 4184
rect 6090 4174 6102 4176
rect 6122 4244 6134 4246
rect 6122 4236 6124 4244
rect 6132 4236 6134 4244
rect 6122 4144 6134 4236
rect 6122 4136 6124 4144
rect 6132 4136 6134 4144
rect 6122 4134 6134 4136
rect 6058 3576 6060 3584
rect 6068 3576 6070 3584
rect 6058 3574 6070 3576
rect 6090 4104 6102 4106
rect 6090 4096 6092 4104
rect 6100 4096 6102 4104
rect 6026 3216 6028 3224
rect 6036 3216 6038 3224
rect 6026 3214 6038 3216
rect 6058 3544 6070 3546
rect 6058 3536 6060 3544
rect 6068 3536 6070 3544
rect 6058 3204 6070 3536
rect 6058 3196 6060 3204
rect 6068 3196 6070 3204
rect 6058 3194 6070 3196
rect 5994 3156 5996 3164
rect 6004 3156 6006 3164
rect 5994 3154 6006 3156
rect 6058 3144 6070 3146
rect 6058 3136 6060 3144
rect 6068 3136 6070 3144
rect 5962 3036 5964 3044
rect 5972 3036 5974 3044
rect 5962 3034 5974 3036
rect 5994 3124 6006 3126
rect 5994 3116 5996 3124
rect 6004 3116 6006 3124
rect 5930 2984 5942 2986
rect 5930 2976 5932 2984
rect 5940 2976 5942 2984
rect 5930 2904 5942 2976
rect 5930 2896 5932 2904
rect 5940 2896 5942 2904
rect 5930 2894 5942 2896
rect 5962 2944 5974 2946
rect 5962 2936 5964 2944
rect 5972 2936 5974 2944
rect 5898 2716 5900 2724
rect 5908 2716 5910 2724
rect 5898 2714 5910 2716
rect 5930 2664 5942 2666
rect 5930 2656 5932 2664
rect 5940 2656 5942 2664
rect 5898 2624 5910 2626
rect 5898 2616 5900 2624
rect 5908 2616 5910 2624
rect 5898 2384 5910 2616
rect 5898 2376 5900 2384
rect 5908 2376 5910 2384
rect 5898 2374 5910 2376
rect 5898 2324 5910 2326
rect 5898 2316 5900 2324
rect 5908 2316 5910 2324
rect 5898 2244 5910 2316
rect 5930 2324 5942 2656
rect 5930 2316 5932 2324
rect 5940 2316 5942 2324
rect 5930 2314 5942 2316
rect 5962 2484 5974 2936
rect 5994 2924 6006 3116
rect 5994 2916 5996 2924
rect 6004 2916 6006 2924
rect 5994 2914 6006 2916
rect 6026 3124 6038 3126
rect 6026 3116 6028 3124
rect 6036 3116 6038 3124
rect 5994 2764 6006 2766
rect 5994 2756 5996 2764
rect 6004 2756 6006 2764
rect 5994 2704 6006 2756
rect 5994 2696 5996 2704
rect 6004 2696 6006 2704
rect 5994 2694 6006 2696
rect 5962 2476 5964 2484
rect 5972 2476 5974 2484
rect 5898 2236 5900 2244
rect 5908 2236 5910 2244
rect 5898 2234 5910 2236
rect 5962 2224 5974 2476
rect 5994 2584 6006 2586
rect 5994 2576 5996 2584
rect 6004 2576 6006 2584
rect 5994 2304 6006 2576
rect 6026 2564 6038 3116
rect 6058 2924 6070 3136
rect 6090 2964 6102 4096
rect 6122 4104 6134 4106
rect 6122 4096 6124 4104
rect 6132 4096 6134 4104
rect 6122 3924 6134 4096
rect 6122 3916 6124 3924
rect 6132 3916 6134 3924
rect 6122 3914 6134 3916
rect 6122 3884 6134 3886
rect 6122 3876 6124 3884
rect 6132 3876 6134 3884
rect 6122 3684 6134 3876
rect 6122 3676 6124 3684
rect 6132 3676 6134 3684
rect 6122 3674 6134 3676
rect 6122 3544 6134 3546
rect 6122 3536 6124 3544
rect 6132 3536 6134 3544
rect 6122 3424 6134 3536
rect 6122 3416 6124 3424
rect 6132 3416 6134 3424
rect 6122 3414 6134 3416
rect 6090 2956 6092 2964
rect 6100 2956 6102 2964
rect 6090 2954 6102 2956
rect 6122 3364 6134 3366
rect 6122 3356 6124 3364
rect 6132 3356 6134 3364
rect 6058 2916 6060 2924
rect 6068 2916 6070 2924
rect 6058 2914 6070 2916
rect 6122 2864 6134 3356
rect 6154 3224 6166 4536
rect 6186 3624 6198 5236
rect 6218 5064 6230 5296
rect 6250 5224 6262 5536
rect 6250 5216 6252 5224
rect 6260 5216 6262 5224
rect 6250 5214 6262 5216
rect 6218 5056 6220 5064
rect 6228 5056 6230 5064
rect 6218 5054 6230 5056
rect 6250 5104 6262 5106
rect 6250 5096 6252 5104
rect 6260 5096 6262 5104
rect 6218 4984 6230 4986
rect 6218 4976 6220 4984
rect 6228 4976 6230 4984
rect 6218 4884 6230 4976
rect 6218 4876 6220 4884
rect 6228 4876 6230 4884
rect 6218 4874 6230 4876
rect 6186 3616 6188 3624
rect 6196 3616 6198 3624
rect 6186 3614 6198 3616
rect 6218 4704 6230 4706
rect 6218 4696 6220 4704
rect 6228 4696 6230 4704
rect 6154 3216 6156 3224
rect 6164 3216 6166 3224
rect 6154 3214 6166 3216
rect 6186 3324 6198 3326
rect 6186 3316 6188 3324
rect 6196 3316 6198 3324
rect 6122 2856 6124 2864
rect 6132 2856 6134 2864
rect 6122 2854 6134 2856
rect 6154 2864 6166 2866
rect 6154 2856 6156 2864
rect 6164 2856 6166 2864
rect 6122 2744 6134 2746
rect 6122 2736 6124 2744
rect 6132 2736 6134 2744
rect 6026 2556 6028 2564
rect 6036 2556 6038 2564
rect 6026 2554 6038 2556
rect 6058 2724 6070 2726
rect 6058 2716 6060 2724
rect 6068 2716 6070 2724
rect 6058 2444 6070 2716
rect 6090 2724 6102 2726
rect 6090 2716 6092 2724
rect 6100 2716 6102 2724
rect 6090 2684 6102 2716
rect 6090 2676 6092 2684
rect 6100 2676 6102 2684
rect 6090 2674 6102 2676
rect 6122 2684 6134 2736
rect 6122 2676 6124 2684
rect 6132 2676 6134 2684
rect 6122 2674 6134 2676
rect 6122 2524 6134 2526
rect 6122 2516 6124 2524
rect 6132 2516 6134 2524
rect 6058 2436 6060 2444
rect 6068 2436 6070 2444
rect 6058 2434 6070 2436
rect 6090 2444 6102 2446
rect 6090 2436 6092 2444
rect 6100 2436 6102 2444
rect 6058 2404 6070 2406
rect 6058 2396 6060 2404
rect 6068 2396 6070 2404
rect 5994 2296 5996 2304
rect 6004 2296 6006 2304
rect 5994 2294 6006 2296
rect 6026 2364 6038 2366
rect 6026 2356 6028 2364
rect 6036 2356 6038 2364
rect 5962 2216 5964 2224
rect 5972 2216 5974 2224
rect 5962 2214 5974 2216
rect 6026 2224 6038 2356
rect 6026 2216 6028 2224
rect 6036 2216 6038 2224
rect 6026 2214 6038 2216
rect 5994 2144 6006 2146
rect 5994 2136 5996 2144
rect 6004 2136 6006 2144
rect 5962 2104 5974 2106
rect 5962 2096 5964 2104
rect 5972 2096 5974 2104
rect 5930 2004 5942 2006
rect 5930 1996 5932 2004
rect 5940 1996 5942 2004
rect 5930 1904 5942 1996
rect 5930 1896 5932 1904
rect 5940 1896 5942 1904
rect 5930 1894 5942 1896
rect 5866 1676 5868 1684
rect 5876 1676 5878 1684
rect 5866 1674 5878 1676
rect 5898 1864 5910 1866
rect 5898 1856 5900 1864
rect 5908 1856 5910 1864
rect 5898 1624 5910 1856
rect 5898 1616 5900 1624
rect 5908 1616 5910 1624
rect 5898 1614 5910 1616
rect 5930 1804 5942 1806
rect 5930 1796 5932 1804
rect 5940 1796 5942 1804
rect 5898 1584 5910 1586
rect 5898 1576 5900 1584
rect 5908 1576 5910 1584
rect 5834 296 5836 304
rect 5844 296 5846 304
rect 5834 294 5846 296
rect 5866 1524 5878 1526
rect 5866 1516 5868 1524
rect 5876 1516 5878 1524
rect 5802 116 5804 124
rect 5812 116 5814 124
rect 5802 114 5814 116
rect 5642 96 5644 104
rect 5652 96 5654 104
rect 5642 94 5654 96
rect 5866 104 5878 1516
rect 5898 624 5910 1576
rect 5898 616 5900 624
rect 5908 616 5910 624
rect 5898 614 5910 616
rect 5898 404 5910 406
rect 5898 396 5900 404
rect 5908 396 5910 404
rect 5898 164 5910 396
rect 5930 404 5942 1796
rect 5962 744 5974 2096
rect 5994 1844 6006 2136
rect 6026 2004 6038 2006
rect 6026 1996 6028 2004
rect 6036 1996 6038 2004
rect 6026 1884 6038 1996
rect 6026 1876 6028 1884
rect 6036 1876 6038 1884
rect 6026 1874 6038 1876
rect 5994 1836 5996 1844
rect 6004 1836 6006 1844
rect 5994 1834 6006 1836
rect 5962 736 5964 744
rect 5972 736 5974 744
rect 5962 734 5974 736
rect 5994 1504 6006 1506
rect 5994 1496 5996 1504
rect 6004 1496 6006 1504
rect 5930 396 5932 404
rect 5940 396 5942 404
rect 5930 394 5942 396
rect 5962 584 5974 586
rect 5962 576 5964 584
rect 5972 576 5974 584
rect 5898 156 5900 164
rect 5908 156 5910 164
rect 5898 154 5910 156
rect 5866 96 5868 104
rect 5876 96 5878 104
rect 5866 94 5878 96
rect 4810 16 4812 24
rect 4820 16 4822 24
rect 4810 14 4822 16
rect 5962 24 5974 576
rect 5994 124 6006 1496
rect 6026 1464 6038 1466
rect 6026 1456 6028 1464
rect 6036 1456 6038 1464
rect 6026 164 6038 1456
rect 6058 1424 6070 2396
rect 6090 2244 6102 2436
rect 6122 2444 6134 2516
rect 6154 2504 6166 2856
rect 6186 2644 6198 3316
rect 6186 2636 6188 2644
rect 6196 2636 6198 2644
rect 6186 2634 6198 2636
rect 6218 2924 6230 4696
rect 6250 4264 6262 5096
rect 6250 4256 6252 4264
rect 6260 4256 6262 4264
rect 6250 4254 6262 4256
rect 6250 4164 6262 4166
rect 6250 4156 6252 4164
rect 6260 4156 6262 4164
rect 6250 4104 6262 4156
rect 6250 4096 6252 4104
rect 6260 4096 6262 4104
rect 6250 4094 6262 4096
rect 6250 3944 6262 3946
rect 6250 3936 6252 3944
rect 6260 3936 6262 3944
rect 6250 3784 6262 3936
rect 6250 3776 6252 3784
rect 6260 3776 6262 3784
rect 6250 3774 6262 3776
rect 6250 3744 6262 3746
rect 6250 3736 6252 3744
rect 6260 3736 6262 3744
rect 6250 3604 6262 3736
rect 6250 3596 6252 3604
rect 6260 3596 6262 3604
rect 6250 3594 6262 3596
rect 6218 2916 6220 2924
rect 6228 2916 6230 2924
rect 6154 2496 6156 2504
rect 6164 2496 6166 2504
rect 6154 2494 6166 2496
rect 6186 2524 6198 2526
rect 6186 2516 6188 2524
rect 6196 2516 6198 2524
rect 6122 2436 6124 2444
rect 6132 2436 6134 2444
rect 6122 2434 6134 2436
rect 6154 2364 6166 2366
rect 6154 2356 6156 2364
rect 6164 2356 6166 2364
rect 6154 2264 6166 2356
rect 6154 2256 6156 2264
rect 6164 2256 6166 2264
rect 6154 2254 6166 2256
rect 6090 2236 6092 2244
rect 6100 2236 6102 2244
rect 6090 2234 6102 2236
rect 6090 2204 6102 2206
rect 6090 2196 6092 2204
rect 6100 2196 6102 2204
rect 6090 2124 6102 2196
rect 6154 2204 6166 2206
rect 6154 2196 6156 2204
rect 6164 2196 6166 2204
rect 6090 2116 6092 2124
rect 6100 2116 6102 2124
rect 6090 2114 6102 2116
rect 6122 2124 6134 2126
rect 6122 2116 6124 2124
rect 6132 2116 6134 2124
rect 6058 1416 6060 1424
rect 6068 1416 6070 1424
rect 6058 1414 6070 1416
rect 6090 2044 6102 2046
rect 6090 2036 6092 2044
rect 6100 2036 6102 2044
rect 6090 884 6102 2036
rect 6122 1984 6134 2116
rect 6122 1976 6124 1984
rect 6132 1976 6134 1984
rect 6122 1974 6134 1976
rect 6122 1924 6134 1926
rect 6122 1916 6124 1924
rect 6132 1916 6134 1924
rect 6122 1884 6134 1916
rect 6154 1904 6166 2196
rect 6154 1896 6156 1904
rect 6164 1896 6166 1904
rect 6154 1894 6166 1896
rect 6122 1876 6124 1884
rect 6132 1876 6134 1884
rect 6122 1874 6134 1876
rect 6186 1864 6198 2516
rect 6186 1856 6188 1864
rect 6196 1856 6198 1864
rect 6186 1854 6198 1856
rect 6218 1904 6230 2916
rect 6218 1896 6220 1904
rect 6228 1896 6230 1904
rect 6090 876 6092 884
rect 6100 876 6102 884
rect 6090 874 6102 876
rect 6122 1684 6134 1686
rect 6122 1676 6124 1684
rect 6132 1676 6134 1684
rect 6026 156 6028 164
rect 6036 156 6038 164
rect 6026 154 6038 156
rect 6058 844 6070 846
rect 6058 836 6060 844
rect 6068 836 6070 844
rect 6058 144 6070 836
rect 6122 644 6134 1676
rect 6154 1484 6166 1486
rect 6154 1476 6156 1484
rect 6164 1476 6166 1484
rect 6154 924 6166 1476
rect 6154 916 6156 924
rect 6164 916 6166 924
rect 6154 914 6166 916
rect 6186 1024 6198 1026
rect 6186 1016 6188 1024
rect 6196 1016 6198 1024
rect 6122 636 6124 644
rect 6132 636 6134 644
rect 6122 634 6134 636
rect 6154 824 6166 826
rect 6154 816 6156 824
rect 6164 816 6166 824
rect 6154 524 6166 816
rect 6154 516 6156 524
rect 6164 516 6166 524
rect 6154 514 6166 516
rect 6186 504 6198 1016
rect 6218 724 6230 1896
rect 6218 716 6220 724
rect 6228 716 6230 724
rect 6218 714 6230 716
rect 6250 3484 6262 3486
rect 6250 3476 6252 3484
rect 6260 3476 6262 3484
rect 6186 496 6188 504
rect 6196 496 6198 504
rect 6186 494 6198 496
rect 6250 324 6262 3476
rect 6250 316 6252 324
rect 6260 316 6262 324
rect 6250 314 6262 316
rect 6058 136 6060 144
rect 6068 136 6070 144
rect 6058 134 6070 136
rect 6154 204 6166 206
rect 6154 196 6156 204
rect 6164 196 6166 204
rect 5994 116 5996 124
rect 6004 116 6006 124
rect 5994 114 6006 116
rect 5962 16 5964 24
rect 5972 16 5974 24
rect 5962 14 5974 16
rect 6154 24 6166 196
rect 6154 16 6156 24
rect 6164 16 6166 24
rect 6154 14 6166 16
rect 4632 6 4636 14
rect 4644 6 4652 14
rect 4660 6 4668 14
rect 4676 6 4680 14
rect 4632 -40 4680 6
use NOR3X1  NOR3X1_3
timestamp 1651764895
transform -1 0 136 0 -1 210
box -4 -6 132 206
use OAI21X1  OAI21X1_77
timestamp 1651764895
transform 1 0 136 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_95
timestamp 1651764895
transform -1 0 264 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_46
timestamp 1651764895
transform -1 0 72 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_23
timestamp 1651764895
transform 1 0 72 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_24
timestamp 1651764895
transform 1 0 136 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_50
timestamp 1651764895
transform 1 0 200 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_76
timestamp 1651764895
transform 1 0 264 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_41
timestamp 1651764895
transform -1 0 392 0 -1 210
box -4 -6 68 206
use OR2X2  OR2X2_10
timestamp 1651764895
transform -1 0 456 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_21
timestamp 1651764895
transform -1 0 328 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_20
timestamp 1651764895
transform -1 0 392 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_14
timestamp 1651764895
transform 1 0 392 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_59
timestamp 1651764895
transform 1 0 456 0 -1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_26
timestamp 1651764895
transform 1 0 504 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_51
timestamp 1651764895
transform 1 0 568 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_83
timestamp 1651764895
transform -1 0 520 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_85
timestamp 1651764895
transform -1 0 584 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_57
timestamp 1651764895
transform -1 0 648 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_20
timestamp 1651764895
transform 1 0 632 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1651764895
transform -1 0 760 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_67
timestamp 1651764895
transform -1 0 824 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_57
timestamp 1651764895
transform -1 0 696 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_85
timestamp 1651764895
transform 1 0 696 0 1 210
box -4 -6 52 206
use INVX1  INVX1_98
timestamp 1651764895
transform 1 0 744 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_134
timestamp 1651764895
transform 1 0 776 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_52
timestamp 1651764895
transform -1 0 888 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_55
timestamp 1651764895
transform 1 0 888 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_105
timestamp 1651764895
transform 1 0 952 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_77
timestamp 1651764895
transform 1 0 984 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_97
timestamp 1651764895
transform -1 0 872 0 1 210
box -4 -6 36 206
use INVX1  INVX1_76
timestamp 1651764895
transform 1 0 872 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_51
timestamp 1651764895
transform 1 0 904 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_50
timestamp 1651764895
transform 1 0 968 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_25
timestamp 1651764895
transform 1 0 1016 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_104
timestamp 1651764895
transform -1 0 1112 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_78
timestamp 1651764895
transform -1 0 1176 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_79
timestamp 1651764895
transform 1 0 1176 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_23
timestamp 1651764895
transform 1 0 1032 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_24
timestamp 1651764895
transform -1 0 1160 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_37
timestamp 1651764895
transform -1 0 1224 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_36
timestamp 1651764895
transform 1 0 1240 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_88
timestamp 1651764895
transform 1 0 1304 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_152
timestamp 1651764895
transform 1 0 1352 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_79
timestamp 1651764895
transform 1 0 1400 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_36
timestamp 1651764895
transform 1 0 1224 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_22
timestamp 1651764895
transform -1 0 1352 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_38
timestamp 1651764895
transform -1 0 1416 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_59
timestamp 1651764895
transform 1 0 1480 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_53
timestamp 1651764895
transform 1 0 1416 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_122
timestamp 1651764895
transform 1 0 1448 0 -1 210
box -4 -6 52 206
use FILL  FILL_1_0_0
timestamp 1651764895
transform 1 0 1544 0 1 210
box -4 -6 20 206
use INVX1  INVX1_131
timestamp 1651764895
transform -1 0 1576 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_80
timestamp 1651764895
transform 1 0 1496 0 -1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_56
timestamp 1651764895
transform 1 0 1592 0 1 210
box -4 -6 68 206
use FILL  FILL_1_0_2
timestamp 1651764895
transform 1 0 1576 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1651764895
transform 1 0 1560 0 1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1651764895
transform 1 0 1608 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1651764895
transform 1 0 1592 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_0
timestamp 1651764895
transform 1 0 1576 0 -1 210
box -4 -6 20 206
use XNOR2X1  XNOR2X1_18
timestamp 1651764895
transform 1 0 1624 0 -1 210
box -4 -6 116 206
use XOR2X1  XOR2X1_8
timestamp 1651764895
transform 1 0 1736 0 -1 210
box -4 -6 116 206
use NAND3X1  NAND3X1_58
timestamp 1651764895
transform -1 0 1720 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_89
timestamp 1651764895
transform 1 0 1720 0 1 210
box -4 -6 52 206
use INVX1  INVX1_158
timestamp 1651764895
transform -1 0 1800 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_155
timestamp 1651764895
transform -1 0 1864 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_112
timestamp 1651764895
transform -1 0 1912 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_107
timestamp 1651764895
transform 1 0 1912 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_95
timestamp 1651764895
transform -1 0 1992 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_62
timestamp 1651764895
transform -1 0 2040 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_157
timestamp 1651764895
transform 1 0 1864 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_197
timestamp 1651764895
transform -1 0 1960 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_22
timestamp 1651764895
transform -1 0 2072 0 1 210
box -4 -6 116 206
use NOR2X1  NOR2X1_63
timestamp 1651764895
transform -1 0 2088 0 -1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_16
timestamp 1651764895
transform 1 0 2088 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_106
timestamp 1651764895
transform -1 0 2232 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_130
timestamp 1651764895
transform -1 0 2104 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_134
timestamp 1651764895
transform 1 0 2104 0 1 210
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1651764895
transform 1 0 2152 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_2
timestamp 1651764895
transform 1 0 2184 0 1 210
box -4 -6 52 206
use XOR2X1  XOR2X1_7
timestamp 1651764895
transform 1 0 2232 0 -1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_106
timestamp 1651764895
transform -1 0 2392 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_14
timestamp 1651764895
transform -1 0 2424 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_4
timestamp 1651764895
transform 1 0 2232 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_3
timestamp 1651764895
transform 1 0 2280 0 1 210
box -4 -6 52 206
use INVX1  INVX1_5
timestamp 1651764895
transform 1 0 2328 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_4
timestamp 1651764895
transform 1 0 2360 0 1 210
box -4 -6 68 206
use AND2X2  AND2X2_3
timestamp 1651764895
transform 1 0 2424 0 -1 210
box -4 -6 68 206
use AND2X2  AND2X2_2
timestamp 1651764895
transform -1 0 2552 0 -1 210
box -4 -6 68 206
use OR2X2  OR2X2_2
timestamp 1651764895
transform -1 0 2616 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_2
timestamp 1651764895
transform -1 0 2472 0 1 210
box -4 -6 52 206
use OR2X2  OR2X2_1
timestamp 1651764895
transform 1 0 2472 0 1 210
box -4 -6 68 206
use AND2X2  AND2X2_1
timestamp 1651764895
transform 1 0 2536 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_8
timestamp 1651764895
transform 1 0 2600 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_6
timestamp 1651764895
transform 1 0 2616 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_10
timestamp 1651764895
transform -1 0 2712 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_9
timestamp 1651764895
transform -1 0 2760 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_10
timestamp 1651764895
transform -1 0 2824 0 -1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_1
timestamp 1651764895
transform -1 0 2760 0 1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_7
timestamp 1651764895
transform -1 0 2808 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_11
timestamp 1651764895
transform -1 0 2856 0 1 210
box -4 -6 52 206
use INVX1  INVX1_12
timestamp 1651764895
transform -1 0 2856 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_8
timestamp 1651764895
transform 1 0 2856 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_13
timestamp 1651764895
transform -1 0 2936 0 -1 210
box -4 -6 36 206
use INVX1  INVX1_185
timestamp 1651764895
transform -1 0 2968 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_98
timestamp 1651764895
transform -1 0 3016 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_5
timestamp 1651764895
transform -1 0 2920 0 1 210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_29
timestamp 1651764895
transform -1 0 3032 0 1 210
box -4 -6 116 206
use INVX1  INVX1_186
timestamp 1651764895
transform 1 0 3080 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_99
timestamp 1651764895
transform 1 0 3032 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_82
timestamp 1651764895
transform -1 0 3128 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_189
timestamp 1651764895
transform 1 0 3016 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_244
timestamp 1651764895
transform 1 0 3160 0 1 210
box -4 -6 68 206
use FILL  FILL_1_1_2
timestamp 1651764895
transform 1 0 3144 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1651764895
transform 1 0 3128 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_0
timestamp 1651764895
transform 1 0 3112 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1651764895
transform -1 0 3176 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1651764895
transform -1 0 3160 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_0
timestamp 1651764895
transform -1 0 3144 0 -1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_50
timestamp 1651764895
transform -1 0 3224 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_72
timestamp 1651764895
transform 1 0 3224 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_81
timestamp 1651764895
transform 1 0 3272 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_51
timestamp 1651764895
transform 1 0 3304 0 -1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_13
timestamp 1651764895
transform 1 0 3352 0 -1 210
box -4 -6 116 206
use XOR2X1  XOR2X1_15
timestamp 1651764895
transform -1 0 3336 0 1 210
box -4 -6 116 206
use NAND2X1  NAND2X1_275
timestamp 1651764895
transform 1 0 3336 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_33
timestamp 1651764895
transform 1 0 3384 0 1 210
box -4 -6 116 206
use INVX1  INVX1_80
timestamp 1651764895
transform -1 0 3496 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_246
timestamp 1651764895
transform 1 0 3496 0 -1 210
box -4 -6 52 206
use XOR2X1  XOR2X1_6
timestamp 1651764895
transform 1 0 3544 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_3
timestamp 1651764895
transform 1 0 3496 0 1 210
box -4 -6 36 206
use INVX1  INVX1_219
timestamp 1651764895
transform 1 0 3528 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_109
timestamp 1651764895
transform -1 0 3608 0 1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_108
timestamp 1651764895
transform -1 0 3656 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_82
timestamp 1651764895
transform -1 0 3704 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_37
timestamp 1651764895
transform -1 0 3752 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_48
timestamp 1651764895
transform 1 0 3752 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_56
timestamp 1651764895
transform -1 0 3864 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_298
timestamp 1651764895
transform -1 0 3720 0 1 210
box -4 -6 68 206
use INVX1  INVX1_218
timestamp 1651764895
transform -1 0 3752 0 1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_5
timestamp 1651764895
transform 1 0 3752 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_3
timestamp 1651764895
transform 1 0 3800 0 1 210
box -4 -6 52 206
use INVX1  INVX1_56
timestamp 1651764895
transform 1 0 3864 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_38
timestamp 1651764895
transform -1 0 3944 0 -1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_12
timestamp 1651764895
transform 1 0 3944 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_6
timestamp 1651764895
transform 1 0 3848 0 1 210
box -4 -6 36 206
use INVX1  INVX1_82
timestamp 1651764895
transform -1 0 3912 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_28
timestamp 1651764895
transform -1 0 3976 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_17
timestamp 1651764895
transform 1 0 3976 0 1 210
box -4 -6 68 206
use INVX1  INVX1_55
timestamp 1651764895
transform -1 0 4088 0 -1 210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_7
timestamp 1651764895
transform 1 0 4088 0 -1 210
box -4 -6 116 206
use INVX1  INVX1_32
timestamp 1651764895
transform 1 0 4200 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_39
timestamp 1651764895
transform -1 0 4104 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_59
timestamp 1651764895
transform -1 0 4152 0 1 210
box -4 -6 52 206
use XOR2X1  XOR2X1_5
timestamp 1651764895
transform 1 0 4152 0 1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_29
timestamp 1651764895
transform 1 0 4232 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_28
timestamp 1651764895
transform 1 0 4296 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_33
timestamp 1651764895
transform -1 0 4376 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_27
timestamp 1651764895
transform 1 0 4376 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_57
timestamp 1651764895
transform 1 0 4264 0 1 210
box -4 -6 36 206
use INVX1  INVX1_83
timestamp 1651764895
transform 1 0 4296 0 1 210
box -4 -6 36 206
use NAND3X1  NAND3X1_29
timestamp 1651764895
transform -1 0 4392 0 1 210
box -4 -6 68 206
use INVX1  INVX1_69
timestamp 1651764895
transform -1 0 4424 0 1 210
box -4 -6 36 206
use INVX1  INVX1_84
timestamp 1651764895
transform 1 0 4488 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_61
timestamp 1651764895
transform 1 0 4424 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_18
timestamp 1651764895
transform 1 0 4472 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_27
timestamp 1651764895
transform -1 0 4472 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_6
timestamp 1651764895
transform 1 0 4584 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_57
timestamp 1651764895
transform 1 0 4520 0 1 210
box -4 -6 68 206
use FILL  FILL_0_2_2
timestamp 1651764895
transform -1 0 4616 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_1
timestamp 1651764895
transform -1 0 4600 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_2_0
timestamp 1651764895
transform -1 0 4584 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_19
timestamp 1651764895
transform 1 0 4520 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_2
timestamp 1651764895
transform -1 0 4808 0 -1 210
box -4 -6 196 206
use NOR2X1  NOR2X1_13
timestamp 1651764895
transform -1 0 4856 0 -1 210
box -4 -6 52 206
use FILL  FILL_1_2_0
timestamp 1651764895
transform -1 0 4648 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_1
timestamp 1651764895
transform -1 0 4664 0 1 210
box -4 -6 20 206
use FILL  FILL_1_2_2
timestamp 1651764895
transform -1 0 4680 0 1 210
box -4 -6 20 206
use DFFPOSX1  DFFPOSX1_1
timestamp 1651764895
transform -1 0 4872 0 1 210
box -4 -6 196 206
use INVX1  INVX1_111
timestamp 1651764895
transform 1 0 4856 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_64
timestamp 1651764895
transform -1 0 4936 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_98
timestamp 1651764895
transform -1 0 4984 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_84
timestamp 1651764895
transform 1 0 4984 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_12
timestamp 1651764895
transform -1 0 4920 0 1 210
box -4 -6 52 206
use AND2X2  AND2X2_4
timestamp 1651764895
transform 1 0 4920 0 1 210
box -4 -6 68 206
use INVX1  INVX1_93
timestamp 1651764895
transform -1 0 5016 0 1 210
box -4 -6 36 206
use AOI21X1  AOI21X1_51
timestamp 1651764895
transform -1 0 5080 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_99
timestamp 1651764895
transform 1 0 5048 0 -1 210
box -4 -6 52 206
use AOI21X1  AOI21X1_30
timestamp 1651764895
transform 1 0 5096 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_90
timestamp 1651764895
transform 1 0 5160 0 -1 210
box -4 -6 36 206
use NOR2X1  NOR2X1_65
timestamp 1651764895
transform 1 0 5192 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_87
timestamp 1651764895
transform 1 0 5080 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_120
timestamp 1651764895
transform -1 0 5208 0 1 210
box -4 -6 68 206
use NOR3X1  NOR3X1_10
timestamp 1651764895
transform 1 0 5208 0 1 210
box -4 -6 132 206
use OR2X2  OR2X2_12
timestamp 1651764895
transform 1 0 5240 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_113
timestamp 1651764895
transform 1 0 5304 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_121
timestamp 1651764895
transform -1 0 5400 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_67
timestamp 1651764895
transform -1 0 5464 0 -1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_53
timestamp 1651764895
transform 1 0 5336 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_111
timestamp 1651764895
transform 1 0 5400 0 1 210
box -4 -6 68 206
use INVX1  INVX1_112
timestamp 1651764895
transform -1 0 5496 0 -1 210
box -4 -6 36 206
use AOI22X1  AOI22X1_16
timestamp 1651764895
transform 1 0 5496 0 -1 210
box -4 -6 84 206
use NAND3X1  NAND3X1_113
timestamp 1651764895
transform -1 0 5640 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_66
timestamp 1651764895
transform 1 0 5464 0 1 210
box -4 -6 52 206
use NAND3X1  NAND3X1_112
timestamp 1651764895
transform 1 0 5512 0 1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_122
timestamp 1651764895
transform -1 0 5640 0 1 210
box -4 -6 68 206
use NOR3X1  NOR3X1_12
timestamp 1651764895
transform 1 0 5640 0 -1 210
box -4 -6 132 206
use NOR2X1  NOR2X1_81
timestamp 1651764895
transform -1 0 5816 0 -1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_19
timestamp 1651764895
transform 1 0 5816 0 -1 210
box -4 -6 116 206
use OAI21X1  OAI21X1_85
timestamp 1651764895
transform -1 0 5704 0 1 210
box -4 -6 68 206
use NOR3X1  NOR3X1_11
timestamp 1651764895
transform 1 0 5704 0 1 210
box -4 -6 132 206
use NAND2X1  NAND2X1_197
timestamp 1651764895
transform 1 0 5928 0 -1 210
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_8
timestamp 1651764895
transform 1 0 5976 0 -1 210
box -4 -6 196 206
use OAI21X1  OAI21X1_123
timestamp 1651764895
transform -1 0 5896 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_68
timestamp 1651764895
transform 1 0 5896 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_100
timestamp 1651764895
transform 1 0 5960 0 1 210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_17
timestamp 1651764895
transform -1 0 6120 0 1 210
box -4 -6 116 206
use AOI21X1  AOI21X1_160
timestamp 1651764895
transform 1 0 6168 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_25
timestamp 1651764895
transform 1 0 6120 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_21
timestamp 1651764895
transform 1 0 6168 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_492
timestamp 1651764895
transform -1 0 6264 0 1 210
box -4 -6 52 206
use FILL  FILL_1_1
timestamp 1651764895
transform -1 0 6248 0 -1 210
box -4 -6 20 206
use FILL  FILL_1_2
timestamp 1651764895
transform -1 0 6264 0 -1 210
box -4 -6 20 206
use NOR3X1  NOR3X1_14
timestamp 1651764895
transform -1 0 136 0 -1 610
box -4 -6 132 206
use AOI21X1  AOI21X1_40
timestamp 1651764895
transform -1 0 200 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_49
timestamp 1651764895
transform 1 0 200 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_79
timestamp 1651764895
transform -1 0 328 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_107
timestamp 1651764895
transform -1 0 392 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_106
timestamp 1651764895
transform 1 0 392 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_80
timestamp 1651764895
transform -1 0 520 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_42
timestamp 1651764895
transform 1 0 520 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_82
timestamp 1651764895
transform -1 0 648 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_67
timestamp 1651764895
transform -1 0 712 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_108
timestamp 1651764895
transform -1 0 776 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_109
timestamp 1651764895
transform 1 0 776 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_75
timestamp 1651764895
transform -1 0 904 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_47
timestamp 1651764895
transform 1 0 904 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_89
timestamp 1651764895
transform -1 0 1032 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_86
timestamp 1651764895
transform -1 0 1096 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_88
timestamp 1651764895
transform 1 0 1096 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_156
timestamp 1651764895
transform 1 0 1160 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_68
timestamp 1651764895
transform -1 0 1256 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_84
timestamp 1651764895
transform 1 0 1256 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_92
timestamp 1651764895
transform -1 0 1384 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_87
timestamp 1651764895
transform 1 0 1384 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_27
timestamp 1651764895
transform -1 0 1512 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_68
timestamp 1651764895
transform 1 0 1512 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_0_0
timestamp 1651764895
transform -1 0 1576 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1651764895
transform -1 0 1592 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1651764895
transform -1 0 1608 0 -1 610
box -4 -6 20 206
use INVX1  INVX1_125
timestamp 1651764895
transform -1 0 1640 0 -1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_93
timestamp 1651764895
transform -1 0 1704 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_90
timestamp 1651764895
transform -1 0 1768 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_71
timestamp 1651764895
transform 1 0 1768 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_35
timestamp 1651764895
transform 1 0 1832 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_57
timestamp 1651764895
transform 1 0 1896 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_83
timestamp 1651764895
transform -1 0 2008 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_56
timestamp 1651764895
transform 1 0 2008 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_34
timestamp 1651764895
transform 1 0 2072 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_78
timestamp 1651764895
transform 1 0 2136 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_52
timestamp 1651764895
transform 1 0 2168 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_164
timestamp 1651764895
transform 1 0 2232 0 -1 610
box -4 -6 52 206
use XOR2X1  XOR2X1_10
timestamp 1651764895
transform -1 0 2392 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_70
timestamp 1651764895
transform 1 0 2392 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_135
timestamp 1651764895
transform 1 0 2440 0 -1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_105
timestamp 1651764895
transform -1 0 2552 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_46
timestamp 1651764895
transform 1 0 2552 0 -1 610
box -4 -6 68 206
use XOR2X1  XOR2X1_11
timestamp 1651764895
transform -1 0 2728 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_216
timestamp 1651764895
transform 1 0 2728 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_114
timestamp 1651764895
transform 1 0 2776 0 -1 610
box -4 -6 68 206
use NOR3X1  NOR3X1_6
timestamp 1651764895
transform 1 0 2840 0 -1 610
box -4 -6 132 206
use AND2X2  AND2X2_33
timestamp 1651764895
transform -1 0 3032 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_107
timestamp 1651764895
transform 1 0 3032 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_1_0
timestamp 1651764895
transform -1 0 3096 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1651764895
transform -1 0 3112 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1651764895
transform -1 0 3128 0 -1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_106
timestamp 1651764895
transform -1 0 3192 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_48
timestamp 1651764895
transform 1 0 3192 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_18
timestamp 1651764895
transform 1 0 3256 0 -1 610
box -4 -6 52 206
use XOR2X1  XOR2X1_2
timestamp 1651764895
transform -1 0 3416 0 -1 610
box -4 -6 116 206
use NAND2X1  NAND2X1_20
timestamp 1651764895
transform 1 0 3416 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_19
timestamp 1651764895
transform -1 0 3512 0 -1 610
box -4 -6 52 206
use XOR2X1  XOR2X1_3
timestamp 1651764895
transform 1 0 3512 0 -1 610
box -4 -6 116 206
use NOR3X1  NOR3X1_7
timestamp 1651764895
transform -1 0 3752 0 -1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_116
timestamp 1651764895
transform 1 0 3752 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_128
timestamp 1651764895
transform 1 0 3816 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_47
timestamp 1651764895
transform 1 0 3880 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_107
timestamp 1651764895
transform 1 0 3944 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_27
timestamp 1651764895
transform 1 0 4008 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_73
timestamp 1651764895
transform 1 0 4072 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_74
timestamp 1651764895
transform -1 0 4168 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_66
timestamp 1651764895
transform 1 0 4168 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_26
timestamp 1651764895
transform 1 0 4232 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_64
timestamp 1651764895
transform 1 0 4296 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_49
timestamp 1651764895
transform 1 0 4360 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_108
timestamp 1651764895
transform 1 0 4424 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_115
timestamp 1651764895
transform -1 0 4552 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_96
timestamp 1651764895
transform -1 0 4600 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_97
timestamp 1651764895
transform -1 0 4648 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_2_0
timestamp 1651764895
transform -1 0 4664 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_1
timestamp 1651764895
transform -1 0 4680 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_2_2
timestamp 1651764895
transform -1 0 4696 0 -1 610
box -4 -6 20 206
use INVX1  INVX1_110
timestamp 1651764895
transform -1 0 4728 0 -1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_65
timestamp 1651764895
transform 1 0 4728 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_32
timestamp 1651764895
transform 1 0 4792 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_118
timestamp 1651764895
transform 1 0 4856 0 -1 610
box -4 -6 36 206
use NOR3X1  NOR3X1_8
timestamp 1651764895
transform -1 0 5016 0 -1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_118
timestamp 1651764895
transform 1 0 5016 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_29
timestamp 1651764895
transform -1 0 5144 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_66
timestamp 1651764895
transform 1 0 5144 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_135
timestamp 1651764895
transform 1 0 5208 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_119
timestamp 1651764895
transform 1 0 5240 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_134
timestamp 1651764895
transform 1 0 5304 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_117
timestamp 1651764895
transform 1 0 5336 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_133
timestamp 1651764895
transform 1 0 5400 0 -1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_52
timestamp 1651764895
transform -1 0 5496 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_109
timestamp 1651764895
transform 1 0 5496 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_110
timestamp 1651764895
transform 1 0 5560 0 -1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_54
timestamp 1651764895
transform 1 0 5624 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_92
timestamp 1651764895
transform 1 0 5688 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_124
timestamp 1651764895
transform 1 0 5720 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_86
timestamp 1651764895
transform 1 0 5784 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_52
timestamp 1651764895
transform 1 0 5848 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_89
timestamp 1651764895
transform -1 0 5928 0 -1 610
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_7
timestamp 1651764895
transform 1 0 5928 0 -1 610
box -4 -6 196 206
use BUFX2  BUFX2_24
timestamp 1651764895
transform 1 0 6120 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_27
timestamp 1651764895
transform 1 0 6168 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_427
timestamp 1651764895
transform -1 0 6264 0 -1 610
box -4 -6 52 206
use NOR3X1  NOR3X1_4
timestamp 1651764895
transform -1 0 136 0 1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_74
timestamp 1651764895
transform -1 0 200 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_73
timestamp 1651764895
transform 1 0 200 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_58
timestamp 1651764895
transform 1 0 264 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_81
timestamp 1651764895
transform 1 0 328 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_97
timestamp 1651764895
transform 1 0 392 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_93
timestamp 1651764895
transform -1 0 504 0 1 610
box -4 -6 52 206
use AOI22X1  AOI22X1_9
timestamp 1651764895
transform -1 0 584 0 1 610
box -4 -6 84 206
use NAND2X1  NAND2X1_92
timestamp 1651764895
transform -1 0 632 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_135
timestamp 1651764895
transform 1 0 632 0 1 610
box -4 -6 68 206
use AOI22X1  AOI22X1_14
timestamp 1651764895
transform -1 0 776 0 1 610
box -4 -6 84 206
use NAND2X1  NAND2X1_111
timestamp 1651764895
transform -1 0 824 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_32
timestamp 1651764895
transform 1 0 824 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_67
timestamp 1651764895
transform -1 0 936 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_63
timestamp 1651764895
transform -1 0 984 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_48
timestamp 1651764895
transform -1 0 1048 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_42
timestamp 1651764895
transform 1 0 1048 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_68
timestamp 1651764895
transform -1 0 1176 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_47
timestamp 1651764895
transform -1 0 1224 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_40
timestamp 1651764895
transform -1 0 1288 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_60
timestamp 1651764895
transform 1 0 1288 0 1 610
box -4 -6 52 206
use INVX1  INVX1_47
timestamp 1651764895
transform 1 0 1336 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_13
timestamp 1651764895
transform 1 0 1368 0 1 610
box -4 -6 68 206
use INVX1  INVX1_75
timestamp 1651764895
transform -1 0 1464 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_4
timestamp 1651764895
transform 1 0 1464 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_6
timestamp 1651764895
transform 1 0 1528 0 1 610
box -4 -6 68 206
use FILL  FILL_3_0_0
timestamp 1651764895
transform 1 0 1592 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1651764895
transform 1 0 1608 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1651764895
transform 1 0 1624 0 1 610
box -4 -6 20 206
use INVX1  INVX1_53
timestamp 1651764895
transform 1 0 1640 0 1 610
box -4 -6 36 206
use NOR3X1  NOR3X1_2
timestamp 1651764895
transform 1 0 1672 0 1 610
box -4 -6 132 206
use NAND3X1  NAND3X1_96
timestamp 1651764895
transform -1 0 1864 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_91
timestamp 1651764895
transform -1 0 1928 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_97
timestamp 1651764895
transform 1 0 1928 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_94
timestamp 1651764895
transform -1 0 2056 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_60
timestamp 1651764895
transform 1 0 2056 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_60
timestamp 1651764895
transform 1 0 2120 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_73
timestamp 1651764895
transform -1 0 2216 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_48
timestamp 1651764895
transform -1 0 2264 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_53
timestamp 1651764895
transform 1 0 2264 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_71
timestamp 1651764895
transform 1 0 2328 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_69
timestamp 1651764895
transform 1 0 2376 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_103
timestamp 1651764895
transform -1 0 2488 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_45
timestamp 1651764895
transform 1 0 2488 0 1 610
box -4 -6 68 206
use INVX1  INVX1_132
timestamp 1651764895
transform 1 0 2552 0 1 610
box -4 -6 36 206
use NOR3X1  NOR3X1_5
timestamp 1651764895
transform -1 0 2712 0 1 610
box -4 -6 132 206
use OAI21X1  OAI21X1_113
timestamp 1651764895
transform 1 0 2712 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_35
timestamp 1651764895
transform 1 0 2776 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_94
timestamp 1651764895
transform -1 0 2888 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_25
timestamp 1651764895
transform -1 0 2952 0 1 610
box -4 -6 68 206
use AND2X2  AND2X2_25
timestamp 1651764895
transform 1 0 2952 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_61
timestamp 1651764895
transform 1 0 3016 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_80
timestamp 1651764895
transform 1 0 3064 0 1 610
box -4 -6 68 206
use FILL  FILL_3_1_0
timestamp 1651764895
transform -1 0 3144 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1651764895
transform -1 0 3160 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1651764895
transform -1 0 3176 0 1 610
box -4 -6 20 206
use INVX1  INVX1_96
timestamp 1651764895
transform -1 0 3208 0 1 610
box -4 -6 36 206
use AOI21X1  AOI21X1_33
timestamp 1651764895
transform 1 0 3208 0 1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_63
timestamp 1651764895
transform 1 0 3272 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_28
timestamp 1651764895
transform 1 0 3336 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1651764895
transform 1 0 3400 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_3
timestamp 1651764895
transform 1 0 3448 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_14
timestamp 1651764895
transform 1 0 3512 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_71
timestamp 1651764895
transform -1 0 3608 0 1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_105
timestamp 1651764895
transform 1 0 3608 0 1 610
box -4 -6 52 206
use INVX1  INVX1_122
timestamp 1651764895
transform 1 0 3656 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_69
timestamp 1651764895
transform -1 0 3752 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_55
timestamp 1651764895
transform 1 0 3752 0 1 610
box -4 -6 68 206
use INVX1  INVX1_121
timestamp 1651764895
transform 1 0 3816 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_94
timestamp 1651764895
transform 1 0 3848 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_123
timestamp 1651764895
transform -1 0 3960 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_27
timestamp 1651764895
transform 1 0 3960 0 1 610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_11
timestamp 1651764895
transform 1 0 4024 0 1 610
box -4 -6 116 206
use AND2X2  AND2X2_21
timestamp 1651764895
transform 1 0 4136 0 1 610
box -4 -6 68 206
use INVX1  INVX1_109
timestamp 1651764895
transform 1 0 4200 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_83
timestamp 1651764895
transform 1 0 4232 0 1 610
box -4 -6 68 206
use INVX1  INVX1_108
timestamp 1651764895
transform 1 0 4296 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_49
timestamp 1651764895
transform 1 0 4328 0 1 610
box -4 -6 52 206
use OR2X2  OR2X2_7
timestamp 1651764895
transform 1 0 4376 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_50
timestamp 1651764895
transform 1 0 4440 0 1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_50
timestamp 1651764895
transform 1 0 4488 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_18
timestamp 1651764895
transform 1 0 4552 0 1 610
box -4 -6 68 206
use FILL  FILL_3_2_0
timestamp 1651764895
transform 1 0 4616 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_1
timestamp 1651764895
transform 1 0 4632 0 1 610
box -4 -6 20 206
use FILL  FILL_3_2_2
timestamp 1651764895
transform 1 0 4648 0 1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_30
timestamp 1651764895
transform 1 0 4664 0 1 610
box -4 -6 68 206
use INVX1  INVX1_86
timestamp 1651764895
transform 1 0 4728 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_31
timestamp 1651764895
transform -1 0 4824 0 1 610
box -4 -6 68 206
use INVX1  INVX1_38
timestamp 1651764895
transform 1 0 4824 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_59
timestamp 1651764895
transform 1 0 4856 0 1 610
box -4 -6 68 206
use INVX1  INVX1_85
timestamp 1651764895
transform 1 0 4920 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_58
timestamp 1651764895
transform 1 0 4952 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_125
timestamp 1651764895
transform -1 0 5080 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_78
timestamp 1651764895
transform 1 0 5080 0 1 610
box -4 -6 52 206
use NOR3X1  NOR3X1_9
timestamp 1651764895
transform -1 0 5256 0 1 610
box -4 -6 132 206
use NAND2X1  NAND2X1_75
timestamp 1651764895
transform 1 0 5256 0 1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_32
timestamp 1651764895
transform -1 0 5368 0 1 610
box -4 -6 68 206
use INVX1  INVX1_87
timestamp 1651764895
transform 1 0 5368 0 1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_76
timestamp 1651764895
transform 1 0 5400 0 1 610
box -4 -6 52 206
use AOI22X1  AOI22X1_4
timestamp 1651764895
transform 1 0 5448 0 1 610
box -4 -6 84 206
use NAND3X1  NAND3X1_33
timestamp 1651764895
transform 1 0 5528 0 1 610
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_6
timestamp 1651764895
transform 1 0 5592 0 1 610
box -4 -6 196 206
use XNOR2X1  XNOR2X1_14
timestamp 1651764895
transform -1 0 5896 0 1 610
box -4 -6 116 206
use BUFX2  BUFX2_23
timestamp 1651764895
transform 1 0 5896 0 1 610
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_9
timestamp 1651764895
transform 1 0 5944 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_26
timestamp 1651764895
transform 1 0 6136 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_310
timestamp 1651764895
transform 1 0 6184 0 1 610
box -4 -6 68 206
use FILL  FILL_4_1
timestamp 1651764895
transform 1 0 6248 0 1 610
box -4 -6 20 206
use NAND3X1  NAND3X1_45
timestamp 1651764895
transform -1 0 72 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_42
timestamp 1651764895
transform -1 0 136 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_65
timestamp 1651764895
transform -1 0 200 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_78
timestamp 1651764895
transform -1 0 264 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_77
timestamp 1651764895
transform 1 0 264 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_37
timestamp 1651764895
transform 1 0 328 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_48
timestamp 1651764895
transform -1 0 456 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_40
timestamp 1651764895
transform -1 0 520 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_47
timestamp 1651764895
transform 1 0 520 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_39
timestamp 1651764895
transform -1 0 648 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_99
timestamp 1651764895
transform -1 0 680 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_96
timestamp 1651764895
transform -1 0 744 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_15
timestamp 1651764895
transform 1 0 744 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_46
timestamp 1651764895
transform -1 0 856 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_18
timestamp 1651764895
transform -1 0 920 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_72
timestamp 1651764895
transform -1 0 952 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_15
timestamp 1651764895
transform 1 0 952 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_61
timestamp 1651764895
transform 1 0 1016 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_49
timestamp 1651764895
transform 1 0 1064 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_5
timestamp 1651764895
transform -1 0 1160 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_10
timestamp 1651764895
transform -1 0 1224 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_42
timestamp 1651764895
transform 1 0 1224 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_43
timestamp 1651764895
transform -1 0 1320 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_54
timestamp 1651764895
transform 1 0 1320 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_7
timestamp 1651764895
transform -1 0 1416 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_54
timestamp 1651764895
transform 1 0 1416 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_44
timestamp 1651764895
transform -1 0 1512 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_27
timestamp 1651764895
transform -1 0 1576 0 -1 1010
box -4 -6 68 206
use FILL  FILL_4_0_0
timestamp 1651764895
transform 1 0 1576 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1651764895
transform 1 0 1592 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1651764895
transform 1 0 1608 0 -1 1010
box -4 -6 20 206
use NAND2X1  NAND2X1_44
timestamp 1651764895
transform 1 0 1624 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_45
timestamp 1651764895
transform -1 0 1720 0 -1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_15
timestamp 1651764895
transform 1 0 1720 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_8
timestamp 1651764895
transform 1 0 1784 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_98
timestamp 1651764895
transform -1 0 1912 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_100
timestamp 1651764895
transform -1 0 1976 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_72
timestamp 1651764895
transform 1 0 1976 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_46
timestamp 1651764895
transform 1 0 2040 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_13
timestamp 1651764895
transform 1 0 2088 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_61
timestamp 1651764895
transform -1 0 2216 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_110
timestamp 1651764895
transform -1 0 2280 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_111
timestamp 1651764895
transform 1 0 2280 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_102
timestamp 1651764895
transform -1 0 2408 0 -1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_15
timestamp 1651764895
transform -1 0 2488 0 -1 1010
box -4 -6 84 206
use INVX1  INVX1_123
timestamp 1651764895
transform -1 0 2520 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_104
timestamp 1651764895
transform 1 0 2520 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_72
timestamp 1651764895
transform -1 0 2632 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_81
timestamp 1651764895
transform 1 0 2632 0 -1 1010
box -4 -6 68 206
use OR2X2  OR2X2_11
timestamp 1651764895
transform 1 0 2696 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_62
timestamp 1651764895
transform -1 0 2824 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_56
timestamp 1651764895
transform -1 0 2872 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_9
timestamp 1651764895
transform 1 0 2872 0 -1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_1
timestamp 1651764895
transform -1 0 3032 0 -1 1010
box -4 -6 116 206
use INVX1  INVX1_25
timestamp 1651764895
transform 1 0 3032 0 -1 1010
box -4 -6 36 206
use FILL  FILL_4_1_0
timestamp 1651764895
transform 1 0 3064 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1651764895
transform 1 0 3080 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1651764895
transform 1 0 3096 0 -1 1010
box -4 -6 20 206
use XNOR2X1  XNOR2X1_3
timestamp 1651764895
transform 1 0 3112 0 -1 1010
box -4 -6 116 206
use OAI21X1  OAI21X1_13
timestamp 1651764895
transform 1 0 3224 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1651764895
transform 1 0 3288 0 -1 1010
box -4 -6 52 206
use OR2X2  OR2X2_4
timestamp 1651764895
transform -1 0 3400 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_15
timestamp 1651764895
transform -1 0 3448 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_55
timestamp 1651764895
transform 1 0 3448 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_49
timestamp 1651764895
transform -1 0 3560 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_54
timestamp 1651764895
transform 1 0 3560 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_70
timestamp 1651764895
transform -1 0 3656 0 -1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_19
timestamp 1651764895
transform 1 0 3656 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_79
timestamp 1651764895
transform 1 0 3720 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_26
timestamp 1651764895
transform -1 0 3816 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_119
timestamp 1651764895
transform 1 0 3816 0 -1 1010
box -4 -6 36 206
use OR2X2  OR2X2_9
timestamp 1651764895
transform 1 0 3848 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_81
timestamp 1651764895
transform 1 0 3912 0 -1 1010
box -4 -6 52 206
use NAND3X1  NAND3X1_34
timestamp 1651764895
transform -1 0 4024 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_31
timestamp 1651764895
transform 1 0 4024 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_55
timestamp 1651764895
transform -1 0 4136 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_65
timestamp 1651764895
transform 1 0 4136 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_94
timestamp 1651764895
transform -1 0 4232 0 -1 1010
box -4 -6 36 206
use XNOR2X1  XNOR2X1_8
timestamp 1651764895
transform 1 0 4232 0 -1 1010
box -4 -6 116 206
use NAND2X1  NAND2X1_35
timestamp 1651764895
transform -1 0 4392 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_40
timestamp 1651764895
transform 1 0 4392 0 -1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_39
timestamp 1651764895
transform 1 0 4424 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_51
timestamp 1651764895
transform 1 0 4472 0 -1 1010
box -4 -6 52 206
use AOI21X1  AOI21X1_9
timestamp 1651764895
transform -1 0 4584 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_64
timestamp 1651764895
transform 1 0 4584 0 -1 1010
box -4 -6 36 206
use INVX1  INVX1_58
timestamp 1651764895
transform 1 0 4616 0 -1 1010
box -4 -6 36 206
use FILL  FILL_4_2_0
timestamp 1651764895
transform 1 0 4648 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_1
timestamp 1651764895
transform 1 0 4664 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_2_2
timestamp 1651764895
transform 1 0 4680 0 -1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_40
timestamp 1651764895
transform 1 0 4696 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_30
timestamp 1651764895
transform 1 0 4744 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_39
timestamp 1651764895
transform -1 0 4840 0 -1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_34
timestamp 1651764895
transform -1 0 4888 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_52
timestamp 1651764895
transform 1 0 4888 0 -1 1010
box -4 -6 52 206
use AND2X2  AND2X2_14
timestamp 1651764895
transform 1 0 4936 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_7
timestamp 1651764895
transform 1 0 5000 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_9
timestamp 1651764895
transform -1 0 5128 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_34
timestamp 1651764895
transform 1 0 5128 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_31
timestamp 1651764895
transform 1 0 5192 0 -1 1010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_9
timestamp 1651764895
transform -1 0 5352 0 -1 1010
box -4 -6 116 206
use OAI21X1  OAI21X1_32
timestamp 1651764895
transform -1 0 5416 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_42
timestamp 1651764895
transform 1 0 5416 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_21
timestamp 1651764895
transform -1 0 5512 0 -1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_17
timestamp 1651764895
transform 1 0 5512 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_88
timestamp 1651764895
transform -1 0 5592 0 -1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_12
timestamp 1651764895
transform -1 0 5656 0 -1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_8
timestamp 1651764895
transform 1 0 5656 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_41
timestamp 1651764895
transform 1 0 5720 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_63
timestamp 1651764895
transform -1 0 5800 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_5
timestamp 1651764895
transform 1 0 5800 0 -1 1010
box -4 -6 196 206
use XNOR2X1  XNOR2X1_23
timestamp 1651764895
transform -1 0 6104 0 -1 1010
box -4 -6 116 206
use BUFX2  BUFX2_22
timestamp 1651764895
transform 1 0 6104 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_129
timestamp 1651764895
transform 1 0 6152 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_20
timestamp 1651764895
transform 1 0 6200 0 -1 1010
box -4 -6 52 206
use FILL  FILL_5_1
timestamp 1651764895
transform -1 0 6264 0 -1 1010
box -4 -6 20 206
use NOR3X1  NOR3X1_13
timestamp 1651764895
transform -1 0 136 0 1 1010
box -4 -6 132 206
use OAI21X1  OAI21X1_103
timestamp 1651764895
transform 1 0 136 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_105
timestamp 1651764895
transform 1 0 200 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_13
timestamp 1651764895
transform -1 0 344 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_120
timestamp 1651764895
transform -1 0 392 0 1 1010
box -4 -6 52 206
use AOI22X1  AOI22X1_12
timestamp 1651764895
transform -1 0 472 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_119
timestamp 1651764895
transform 1 0 472 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_22
timestamp 1651764895
transform -1 0 584 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_87
timestamp 1651764895
transform 1 0 584 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_70
timestamp 1651764895
transform -1 0 696 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_69
timestamp 1651764895
transform -1 0 760 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_110
timestamp 1651764895
transform -1 0 808 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_62
timestamp 1651764895
transform -1 0 856 0 1 1010
box -4 -6 52 206
use OAI22X1  OAI22X1_4
timestamp 1651764895
transform 1 0 856 0 1 1010
box -4 -6 84 206
use NAND2X1  NAND2X1_86
timestamp 1651764895
transform -1 0 984 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_41
timestamp 1651764895
transform 1 0 984 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_16
timestamp 1651764895
transform 1 0 1048 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_37
timestamp 1651764895
transform -1 0 1160 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_15
timestamp 1651764895
transform 1 0 1160 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_16
timestamp 1651764895
transform -1 0 1256 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_23
timestamp 1651764895
transform 1 0 1256 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_30
timestamp 1651764895
transform -1 0 1352 0 1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_70
timestamp 1651764895
transform -1 0 1416 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_138
timestamp 1651764895
transform -1 0 1480 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_140
timestamp 1651764895
transform -1 0 1544 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1651764895
transform 1 0 1544 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1651764895
transform 1 0 1560 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1651764895
transform 1 0 1576 0 1 1010
box -4 -6 20 206
use AOI21X1  AOI21X1_69
timestamp 1651764895
transform 1 0 1592 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_153
timestamp 1651764895
transform 1 0 1656 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_154
timestamp 1651764895
transform 1 0 1720 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_144
timestamp 1651764895
transform -1 0 1848 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_141
timestamp 1651764895
transform 1 0 1848 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_145
timestamp 1651764895
transform -1 0 1976 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_148
timestamp 1651764895
transform -1 0 2040 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_142
timestamp 1651764895
transform -1 0 2104 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_143
timestamp 1651764895
transform -1 0 2168 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_149
timestamp 1651764895
transform -1 0 2232 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_151
timestamp 1651764895
transform 1 0 2232 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_146
timestamp 1651764895
transform -1 0 2360 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_99
timestamp 1651764895
transform 1 0 2360 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_95
timestamp 1651764895
transform 1 0 2424 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_43
timestamp 1651764895
transform 1 0 2488 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_159
timestamp 1651764895
transform 1 0 2552 0 1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_74
timestamp 1651764895
transform -1 0 2648 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_160
timestamp 1651764895
transform 1 0 2648 0 1 1010
box -4 -6 68 206
use NOR3X1  NOR3X1_15
timestamp 1651764895
transform -1 0 2840 0 1 1010
box -4 -6 132 206
use OAI21X1  OAI21X1_157
timestamp 1651764895
transform 1 0 2840 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_156
timestamp 1651764895
transform 1 0 2904 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_158
timestamp 1651764895
transform 1 0 2968 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_161
timestamp 1651764895
transform 1 0 3032 0 1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_163
timestamp 1651764895
transform 1 0 3064 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_1_0
timestamp 1651764895
transform -1 0 3144 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1651764895
transform -1 0 3160 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1651764895
transform -1 0 3176 0 1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_161
timestamp 1651764895
transform -1 0 3240 0 1 1010
box -4 -6 68 206
use AOI21X1  AOI21X1_76
timestamp 1651764895
transform 1 0 3240 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_162
timestamp 1651764895
transform 1 0 3304 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_133
timestamp 1651764895
transform -1 0 3416 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_11
timestamp 1651764895
transform 1 0 3416 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1651764895
transform 1 0 3480 0 1 1010
box -4 -6 52 206
use AND2X2  AND2X2_39
timestamp 1651764895
transform 1 0 3528 0 1 1010
box -4 -6 68 206
use AOI22X1  AOI22X1_22
timestamp 1651764895
transform 1 0 3592 0 1 1010
box -4 -6 84 206
use NAND3X1  NAND3X1_164
timestamp 1651764895
transform -1 0 3736 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_160
timestamp 1651764895
transform 1 0 3736 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_163
timestamp 1651764895
transform -1 0 3832 0 1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_16
timestamp 1651764895
transform 1 0 3832 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_44
timestamp 1651764895
transform -1 0 3944 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_47
timestamp 1651764895
transform -1 0 3992 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_68
timestamp 1651764895
transform 1 0 3992 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_28
timestamp 1651764895
transform -1 0 4088 0 1 1010
box -4 -6 68 206
use AND2X2  AND2X2_20
timestamp 1651764895
transform 1 0 4088 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_23
timestamp 1651764895
transform 1 0 4152 0 1 1010
box -4 -6 36 206
use INVX1  INVX1_26
timestamp 1651764895
transform 1 0 4184 0 1 1010
box -4 -6 36 206
use NAND2X1  NAND2X1_23
timestamp 1651764895
transform 1 0 4216 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_31
timestamp 1651764895
transform -1 0 4312 0 1 1010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_5
timestamp 1651764895
transform -1 0 4424 0 1 1010
box -4 -6 116 206
use OAI21X1  OAI21X1_22
timestamp 1651764895
transform -1 0 4488 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_6
timestamp 1651764895
transform 1 0 4488 0 1 1010
box -4 -6 116 206
use NOR2X1  NOR2X1_32
timestamp 1651764895
transform 1 0 4600 0 1 1010
box -4 -6 52 206
use FILL  FILL_5_2_0
timestamp 1651764895
transform -1 0 4664 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_1
timestamp 1651764895
transform -1 0 4680 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_2_2
timestamp 1651764895
transform -1 0 4696 0 1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_33
timestamp 1651764895
transform -1 0 4744 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_28
timestamp 1651764895
transform 1 0 4744 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_29
timestamp 1651764895
transform 1 0 4792 0 1 1010
box -4 -6 52 206
use OR2X2  OR2X2_5
timestamp 1651764895
transform 1 0 4840 0 1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_33
timestamp 1651764895
transform -1 0 4952 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_34
timestamp 1651764895
transform -1 0 5000 0 1 1010
box -4 -6 52 206
use XOR2X1  XOR2X1_4
timestamp 1651764895
transform 1 0 5000 0 1 1010
box -4 -6 116 206
use INVX1  INVX1_35
timestamp 1651764895
transform -1 0 5144 0 1 1010
box -4 -6 36 206
use INVX1  INVX1_59
timestamp 1651764895
transform 1 0 5144 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_31
timestamp 1651764895
transform 1 0 5176 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_24
timestamp 1651764895
transform -1 0 5272 0 1 1010
box -4 -6 36 206
use AOI21X1  AOI21X1_6
timestamp 1651764895
transform 1 0 5272 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1651764895
transform 1 0 5336 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_62
timestamp 1651764895
transform 1 0 5400 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_33
timestamp 1651764895
transform 1 0 5432 0 1 1010
box -4 -6 68 206
use INVX1  INVX1_60
timestamp 1651764895
transform -1 0 5528 0 1 1010
box -4 -6 36 206
use INVX1  INVX1_61
timestamp 1651764895
transform 1 0 5528 0 1 1010
box -4 -6 36 206
use NAND3X1  NAND3X1_11
timestamp 1651764895
transform 1 0 5560 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_29
timestamp 1651764895
transform 1 0 5624 0 1 1010
box -4 -6 52 206
use INVX1  INVX1_21
timestamp 1651764895
transform 1 0 5672 0 1 1010
box -4 -6 36 206
use NOR2X1  NOR2X1_22
timestamp 1651764895
transform 1 0 5704 0 1 1010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_10
timestamp 1651764895
transform -1 0 5864 0 1 1010
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_3
timestamp 1651764895
transform 1 0 5864 0 1 1010
box -4 -6 196 206
use DFFPOSX1  DFFPOSX1_4
timestamp 1651764895
transform 1 0 6056 0 1 1010
box -4 -6 196 206
use FILL  FILL_6_1
timestamp 1651764895
transform 1 0 6248 0 1 1010
box -4 -6 20 206
use INVX1  INVX1_100
timestamp 1651764895
transform 1 0 8 0 -1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_38
timestamp 1651764895
transform 1 0 40 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_41
timestamp 1651764895
transform 1 0 104 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_76
timestamp 1651764895
transform -1 0 232 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_72
timestamp 1651764895
transform 1 0 232 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_141
timestamp 1651764895
transform 1 0 296 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_75
timestamp 1651764895
transform -1 0 424 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_70
timestamp 1651764895
transform -1 0 488 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_99
timestamp 1651764895
transform -1 0 552 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_104
timestamp 1651764895
transform 1 0 552 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_126
timestamp 1651764895
transform 1 0 616 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_112
timestamp 1651764895
transform 1 0 648 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_59
timestamp 1651764895
transform 1 0 696 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_98
timestamp 1651764895
transform -1 0 824 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_46
timestamp 1651764895
transform 1 0 824 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_51
timestamp 1651764895
transform 1 0 888 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_45
timestamp 1651764895
transform -1 0 968 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_49
timestamp 1651764895
transform 1 0 968 0 -1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_1
timestamp 1651764895
transform 1 0 1032 0 -1 1410
box -4 -6 132 206
use NAND3X1  NAND3X1_4
timestamp 1651764895
transform -1 0 1224 0 -1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_2
timestamp 1651764895
transform -1 0 1304 0 -1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_41
timestamp 1651764895
transform -1 0 1352 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_52
timestamp 1651764895
transform -1 0 1384 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_151
timestamp 1651764895
transform -1 0 1448 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_152
timestamp 1651764895
transform 1 0 1448 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_137
timestamp 1651764895
transform -1 0 1576 0 -1 1410
box -4 -6 68 206
use FILL  FILL_6_0_0
timestamp 1651764895
transform -1 0 1592 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1651764895
transform -1 0 1608 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1651764895
transform -1 0 1624 0 -1 1410
box -4 -6 20 206
use NAND3X1  NAND3X1_139
timestamp 1651764895
transform -1 0 1688 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_84
timestamp 1651764895
transform 1 0 1688 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_155
timestamp 1651764895
transform -1 0 1784 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_175
timestamp 1651764895
transform 1 0 1784 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_183
timestamp 1651764895
transform 1 0 1848 0 -1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_95
timestamp 1651764895
transform 1 0 1880 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_2
timestamp 1651764895
transform 1 0 1944 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_16
timestamp 1651764895
transform 1 0 2008 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_25
timestamp 1651764895
transform -1 0 2120 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_17
timestamp 1651764895
transform 1 0 2120 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_83
timestamp 1651764895
transform 1 0 2184 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_9
timestamp 1651764895
transform 1 0 2248 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_18
timestamp 1651764895
transform -1 0 2376 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_31
timestamp 1651764895
transform -1 0 2408 0 -1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_150
timestamp 1651764895
transform -1 0 2472 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_5
timestamp 1651764895
transform -1 0 2536 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_3
timestamp 1651764895
transform 1 0 2536 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_10
timestamp 1651764895
transform 1 0 2600 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_44
timestamp 1651764895
transform -1 0 2728 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_166
timestamp 1651764895
transform 1 0 2728 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_101
timestamp 1651764895
transform -1 0 2840 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_158
timestamp 1651764895
transform 1 0 2840 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_73
timestamp 1651764895
transform 1 0 2904 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_133
timestamp 1651764895
transform 1 0 2968 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_150
timestamp 1651764895
transform -1 0 3080 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_129
timestamp 1651764895
transform 1 0 3080 0 -1 1410
box -4 -6 36 206
use FILL  FILL_6_1_0
timestamp 1651764895
transform 1 0 3112 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1651764895
transform 1 0 3128 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1651764895
transform 1 0 3144 0 -1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_121
timestamp 1651764895
transform 1 0 3160 0 -1 1410
box -4 -6 52 206
use AND2X2  AND2X2_36
timestamp 1651764895
transform 1 0 3208 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_165
timestamp 1651764895
transform 1 0 3272 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_115
timestamp 1651764895
transform -1 0 3384 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_143
timestamp 1651764895
transform -1 0 3416 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_7
timestamp 1651764895
transform -1 0 3464 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_2
timestamp 1651764895
transform 1 0 3464 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_11
timestamp 1651764895
transform 1 0 3528 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_9
timestamp 1651764895
transform -1 0 3624 0 -1 1410
box -4 -6 68 206
use OAI22X1  OAI22X1_1
timestamp 1651764895
transform 1 0 3624 0 -1 1410
box -4 -6 84 206
use OAI22X1  OAI22X1_3
timestamp 1651764895
transform 1 0 3704 0 -1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_160
timestamp 1651764895
transform 1 0 3784 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_165
timestamp 1651764895
transform -1 0 3896 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_75
timestamp 1651764895
transform 1 0 3896 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_67
timestamp 1651764895
transform 1 0 3960 0 -1 1410
box -4 -6 36 206
use AOI22X1  AOI22X1_1
timestamp 1651764895
transform -1 0 4072 0 -1 1410
box -4 -6 84 206
use NOR2X1  NOR2X1_35
timestamp 1651764895
transform 1 0 4072 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_42
timestamp 1651764895
transform -1 0 4152 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_12
timestamp 1651764895
transform 1 0 4152 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_56
timestamp 1651764895
transform 1 0 4216 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_8
timestamp 1651764895
transform 1 0 4264 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_23
timestamp 1651764895
transform -1 0 4376 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_43
timestamp 1651764895
transform 1 0 4376 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_14
timestamp 1651764895
transform 1 0 4424 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_57
timestamp 1651764895
transform 1 0 4488 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_38
timestamp 1651764895
transform 1 0 4536 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_58
timestamp 1651764895
transform -1 0 4648 0 -1 1410
box -4 -6 52 206
use FILL  FILL_6_2_0
timestamp 1651764895
transform 1 0 4648 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_1
timestamp 1651764895
transform 1 0 4664 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_2_2
timestamp 1651764895
transform 1 0 4680 0 -1 1410
box -4 -6 20 206
use AND2X2  AND2X2_19
timestamp 1651764895
transform 1 0 4696 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_30
timestamp 1651764895
transform 1 0 4760 0 -1 1410
box -4 -6 52 206
use OR2X2  OR2X2_6
timestamp 1651764895
transform 1 0 4808 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_11
timestamp 1651764895
transform 1 0 4872 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_34
timestamp 1651764895
transform 1 0 4936 0 -1 1410
box -4 -6 36 206
use AOI21X1  AOI21X1_1
timestamp 1651764895
transform -1 0 5032 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_60
timestamp 1651764895
transform 1 0 5032 0 -1 1410
box -4 -6 68 206
use AND2X2  AND2X2_6
timestamp 1651764895
transform -1 0 5160 0 -1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_53
timestamp 1651764895
transform -1 0 5208 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_101
timestamp 1651764895
transform 1 0 5208 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_69
timestamp 1651764895
transform 1 0 5256 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_102
timestamp 1651764895
transform 1 0 5304 0 -1 1410
box -4 -6 52 206
use NOR3X1  NOR3X1_17
timestamp 1651764895
transform -1 0 5480 0 -1 1410
box -4 -6 132 206
use OAI21X1  OAI21X1_162
timestamp 1651764895
transform 1 0 5480 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_169
timestamp 1651764895
transform -1 0 5608 0 -1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_80
timestamp 1651764895
transform 1 0 5608 0 -1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_19
timestamp 1651764895
transform -1 0 5800 0 -1 1410
box -4 -6 132 206
use OAI21X1  OAI21X1_163
timestamp 1651764895
transform 1 0 5800 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_193
timestamp 1651764895
transform 1 0 5864 0 -1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_81
timestamp 1651764895
transform -1 0 5976 0 -1 1410
box -4 -6 68 206
use INVX1  INVX1_166
timestamp 1651764895
transform -1 0 6008 0 -1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_153
timestamp 1651764895
transform 1 0 6008 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_10
timestamp 1651764895
transform 1 0 6056 0 -1 1410
box -4 -6 196 206
use FILL  FILL_7_1
timestamp 1651764895
transform -1 0 6264 0 -1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_88
timestamp 1651764895
transform -1 0 56 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_72
timestamp 1651764895
transform -1 0 120 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_101
timestamp 1651764895
transform 1 0 120 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_100
timestamp 1651764895
transform 1 0 152 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_22
timestamp 1651764895
transform -1 0 280 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_62
timestamp 1651764895
transform -1 0 344 0 1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_8
timestamp 1651764895
transform -1 0 424 0 1 1410
box -4 -6 84 206
use NAND2X1  NAND2X1_113
timestamp 1651764895
transform -1 0 472 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_77
timestamp 1651764895
transform -1 0 520 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_28
timestamp 1651764895
transform -1 0 584 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_40
timestamp 1651764895
transform -1 0 632 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_23
timestamp 1651764895
transform -1 0 696 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_18
timestamp 1651764895
transform 1 0 696 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_76
timestamp 1651764895
transform 1 0 760 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_109
timestamp 1651764895
transform -1 0 856 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_19
timestamp 1651764895
transform 1 0 856 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_12
timestamp 1651764895
transform -1 0 984 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1651764895
transform 1 0 984 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_24
timestamp 1651764895
transform -1 0 1080 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_24
timestamp 1651764895
transform 1 0 1080 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_25
timestamp 1651764895
transform 1 0 1144 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_26
timestamp 1651764895
transform -1 0 1272 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_15
timestamp 1651764895
transform 1 0 1272 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_3
timestamp 1651764895
transform 1 0 1336 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_48
timestamp 1651764895
transform 1 0 1400 0 1 1410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_4
timestamp 1651764895
transform -1 0 1544 0 1 1410
box -4 -6 116 206
use NOR2X1  NOR2X1_26
timestamp 1651764895
transform -1 0 1592 0 1 1410
box -4 -6 52 206
use FILL  FILL_7_0_0
timestamp 1651764895
transform 1 0 1592 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1651764895
transform 1 0 1608 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1651764895
transform 1 0 1624 0 1 1410
box -4 -6 20 206
use OR2X2  OR2X2_3
timestamp 1651764895
transform 1 0 1640 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_8
timestamp 1651764895
transform 1 0 1704 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_5
timestamp 1651764895
transform 1 0 1768 0 1 1410
box -4 -6 68 206
use AND2X2  AND2X2_7
timestamp 1651764895
transform 1 0 1832 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_36
timestamp 1651764895
transform 1 0 1896 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_24
timestamp 1651764895
transform -1 0 1992 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_8
timestamp 1651764895
transform 1 0 1992 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_17
timestamp 1651764895
transform -1 0 2104 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_12
timestamp 1651764895
transform -1 0 2152 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_15
timestamp 1651764895
transform 1 0 2152 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_18
timestamp 1651764895
transform 1 0 2200 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_17
timestamp 1651764895
transform 1 0 2248 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_154
timestamp 1651764895
transform -1 0 2344 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_147
timestamp 1651764895
transform -1 0 2408 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_152
timestamp 1651764895
transform 1 0 2408 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_142
timestamp 1651764895
transform 1 0 2472 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_151
timestamp 1651764895
transform 1 0 2504 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_149
timestamp 1651764895
transform 1 0 2552 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_159
timestamp 1651764895
transform -1 0 2664 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_160
timestamp 1651764895
transform -1 0 2696 0 1 1410
box -4 -6 36 206
use AOI22X1  AOI22X1_21
timestamp 1651764895
transform -1 0 2776 0 1 1410
box -4 -6 84 206
use NAND3X1  NAND3X1_153
timestamp 1651764895
transform -1 0 2840 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_157
timestamp 1651764895
transform -1 0 2904 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_128
timestamp 1651764895
transform 1 0 2904 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_132
timestamp 1651764895
transform -1 0 3000 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_130
timestamp 1651764895
transform 1 0 3000 0 1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_114
timestamp 1651764895
transform -1 0 3112 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_1_0
timestamp 1651764895
transform -1 0 3128 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1651764895
transform -1 0 3144 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1651764895
transform -1 0 3160 0 1 1410
box -4 -6 20 206
use OAI21X1  OAI21X1_169
timestamp 1651764895
transform -1 0 3224 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_131
timestamp 1651764895
transform 1 0 3224 0 1 1410
box -4 -6 52 206
use AND2X2  AND2X2_35
timestamp 1651764895
transform -1 0 3336 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_129
timestamp 1651764895
transform -1 0 3384 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_26
timestamp 1651764895
transform 1 0 3384 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_80
timestamp 1651764895
transform 1 0 3432 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_129
timestamp 1651764895
transform 1 0 3480 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_104
timestamp 1651764895
transform -1 0 3592 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_93
timestamp 1651764895
transform 1 0 3592 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_54
timestamp 1651764895
transform 1 0 3656 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_95
timestamp 1651764895
transform 1 0 3704 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_90
timestamp 1651764895
transform 1 0 3736 0 1 1410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_15
timestamp 1651764895
transform -1 0 3912 0 1 1410
box -4 -6 116 206
use OAI21X1  OAI21X1_64
timestamp 1651764895
transform 1 0 3912 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_37
timestamp 1651764895
transform 1 0 3976 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_66
timestamp 1651764895
transform 1 0 4040 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_13
timestamp 1651764895
transform -1 0 4136 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_55
timestamp 1651764895
transform 1 0 4136 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_62
timestamp 1651764895
transform -1 0 4248 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1651764895
transform 1 0 4248 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_22
timestamp 1651764895
transform 1 0 4296 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_21
timestamp 1651764895
transform 1 0 4344 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_162
timestamp 1651764895
transform 1 0 4408 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_159
timestamp 1651764895
transform 1 0 4440 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_165
timestamp 1651764895
transform 1 0 4504 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_140
timestamp 1651764895
transform -1 0 4600 0 1 1410
box -4 -6 36 206
use AND2X2  AND2X2_34
timestamp 1651764895
transform -1 0 4664 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_2_0
timestamp 1651764895
transform -1 0 4680 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_1
timestamp 1651764895
transform -1 0 4696 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_2_2
timestamp 1651764895
transform -1 0 4712 0 1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_125
timestamp 1651764895
transform -1 0 4760 0 1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_77
timestamp 1651764895
transform -1 0 4824 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_166
timestamp 1651764895
transform 1 0 4824 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_167
timestamp 1651764895
transform -1 0 4952 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_79
timestamp 1651764895
transform 1 0 4952 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_165
timestamp 1651764895
transform 1 0 5016 0 1 1410
box -4 -6 36 206
use INVX1  INVX1_164
timestamp 1651764895
transform 1 0 5048 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_161
timestamp 1651764895
transform 1 0 5080 0 1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_16
timestamp 1651764895
transform 1 0 5144 0 1 1410
box -4 -6 132 206
use NAND3X1  NAND3X1_168
timestamp 1651764895
transform -1 0 5336 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_78
timestamp 1651764895
transform 1 0 5336 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_117
timestamp 1651764895
transform 1 0 5400 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_164
timestamp 1651764895
transform -1 0 5496 0 1 1410
box -4 -6 68 206
use NOR3X1  NOR3X1_18
timestamp 1651764895
transform -1 0 5624 0 1 1410
box -4 -6 132 206
use INVX1  INVX1_137
timestamp 1651764895
transform -1 0 5656 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_220
timestamp 1651764895
transform -1 0 5720 0 1 1410
box -4 -6 68 206
use AOI21X1  AOI21X1_105
timestamp 1651764895
transform 1 0 5720 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_192
timestamp 1651764895
transform -1 0 5832 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_206
timestamp 1651764895
transform -1 0 5896 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_194
timestamp 1651764895
transform -1 0 5944 0 1 1410
box -4 -6 52 206
use XOR2X1  XOR2X1_12
timestamp 1651764895
transform -1 0 6056 0 1 1410
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_12
timestamp 1651764895
transform 1 0 6056 0 1 1410
box -4 -6 196 206
use FILL  FILL_8_1
timestamp 1651764895
transform 1 0 6248 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_11
timestamp 1651764895
transform 1 0 8 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_13
timestamp 1651764895
transform 1 0 56 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_10
timestamp 1651764895
transform 1 0 104 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_12
timestamp 1651764895
transform 1 0 152 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_44
timestamp 1651764895
transform -1 0 264 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_58
timestamp 1651764895
transform -1 0 312 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_43
timestamp 1651764895
transform 1 0 312 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_1
timestamp 1651764895
transform 1 0 376 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_91
timestamp 1651764895
transform -1 0 456 0 -1 1810
box -4 -6 52 206
use AND2X2  AND2X2_17
timestamp 1651764895
transform 1 0 456 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_103
timestamp 1651764895
transform 1 0 520 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_66
timestamp 1651764895
transform 1 0 552 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_102
timestamp 1651764895
transform 1 0 600 0 -1 1810
box -4 -6 36 206
use AOI22X1  AOI22X1_7
timestamp 1651764895
transform 1 0 632 0 -1 1810
box -4 -6 84 206
use OAI21X1  OAI21X1_71
timestamp 1651764895
transform 1 0 712 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_74
timestamp 1651764895
transform -1 0 808 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_17
timestamp 1651764895
transform 1 0 808 0 -1 1810
box -4 -6 68 206
use AOI22X1  AOI22X1_3
timestamp 1651764895
transform 1 0 872 0 -1 1810
box -4 -6 84 206
use NAND2X1  NAND2X1_64
timestamp 1651764895
transform -1 0 1000 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_44
timestamp 1651764895
transform -1 0 1064 0 -1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_11
timestamp 1651764895
transform -1 0 1128 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_16
timestamp 1651764895
transform 1 0 1128 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_43
timestamp 1651764895
transform -1 0 1256 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_45
timestamp 1651764895
transform -1 0 1320 0 -1 1810
box -4 -6 68 206
use AND2X2  AND2X2_12
timestamp 1651764895
transform -1 0 1384 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_36
timestamp 1651764895
transform -1 0 1432 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_11
timestamp 1651764895
transform 1 0 1432 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_14
timestamp 1651764895
transform 1 0 1480 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_0_0
timestamp 1651764895
transform 1 0 1544 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1651764895
transform 1 0 1560 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1651764895
transform 1 0 1576 0 -1 1810
box -4 -6 20 206
use OAI22X1  OAI22X1_2
timestamp 1651764895
transform 1 0 1592 0 -1 1810
box -4 -6 84 206
use NAND2X1  NAND2X1_5
timestamp 1651764895
transform -1 0 1720 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_4
timestamp 1651764895
transform 1 0 1720 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_7
timestamp 1651764895
transform 1 0 1768 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_6
timestamp 1651764895
transform -1 0 1896 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_1
timestamp 1651764895
transform -1 0 1960 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_16
timestamp 1651764895
transform -1 0 2008 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1651764895
transform -1 0 2072 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_194
timestamp 1651764895
transform -1 0 2136 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_192
timestamp 1651764895
transform -1 0 2200 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_195
timestamp 1651764895
transform -1 0 2264 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_196
timestamp 1651764895
transform 1 0 2264 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_195
timestamp 1651764895
transform -1 0 2392 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_198
timestamp 1651764895
transform 1 0 2392 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_197
timestamp 1651764895
transform 1 0 2456 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_173
timestamp 1651764895
transform 1 0 2520 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_193
timestamp 1651764895
transform -1 0 2616 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_2
timestamp 1651764895
transform 1 0 2616 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_155
timestamp 1651764895
transform -1 0 2744 0 -1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_106
timestamp 1651764895
transform 1 0 2744 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_148
timestamp 1651764895
transform -1 0 2856 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_82
timestamp 1651764895
transform 1 0 2856 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_173
timestamp 1651764895
transform 1 0 2920 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_171
timestamp 1651764895
transform -1 0 3016 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_156
timestamp 1651764895
transform -1 0 3080 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_184
timestamp 1651764895
transform -1 0 3112 0 -1 1810
box -4 -6 36 206
use FILL  FILL_8_1_0
timestamp 1651764895
transform 1 0 3112 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1651764895
transform 1 0 3128 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1651764895
transform 1 0 3144 0 -1 1810
box -4 -6 20 206
use AOI21X1  AOI21X1_100
timestamp 1651764895
transform 1 0 3160 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_167
timestamp 1651764895
transform -1 0 3272 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_187
timestamp 1651764895
transform 1 0 3272 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_198
timestamp 1651764895
transform -1 0 3368 0 -1 1810
box -4 -6 68 206
use NOR3X1  NOR3X1_20
timestamp 1651764895
transform 1 0 3368 0 -1 1810
box -4 -6 132 206
use NOR2X1  NOR2X1_85
timestamp 1651764895
transform 1 0 3496 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_141
timestamp 1651764895
transform 1 0 3544 0 -1 1810
box -4 -6 36 206
use OR2X2  OR2X2_16
timestamp 1651764895
transform -1 0 3640 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_132
timestamp 1651764895
transform -1 0 3704 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_126
timestamp 1651764895
transform -1 0 3752 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_91
timestamp 1651764895
transform 1 0 3752 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_92
timestamp 1651764895
transform -1 0 3880 0 -1 1810
box -4 -6 68 206
use OR2X2  OR2X2_14
timestamp 1651764895
transform -1 0 3944 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_120
timestamp 1651764895
transform -1 0 3976 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_70
timestamp 1651764895
transform -1 0 4024 0 -1 1810
box -4 -6 52 206
use OR2X2  OR2X2_13
timestamp 1651764895
transform -1 0 4088 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_63
timestamp 1651764895
transform -1 0 4152 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_79
timestamp 1651764895
transform -1 0 4200 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_36
timestamp 1651764895
transform 1 0 4200 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_35
timestamp 1651764895
transform -1 0 4328 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_53
timestamp 1651764895
transform -1 0 4376 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_32
timestamp 1651764895
transform 1 0 4376 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_20
timestamp 1651764895
transform -1 0 4488 0 -1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_30
timestamp 1651764895
transform 1 0 4488 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_37
timestamp 1651764895
transform 1 0 4536 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_18
timestamp 1651764895
transform -1 0 4600 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_203
timestamp 1651764895
transform 1 0 4600 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_2_0
timestamp 1651764895
transform -1 0 4680 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_1
timestamp 1651764895
transform -1 0 4696 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_2_2
timestamp 1651764895
transform -1 0 4712 0 -1 1810
box -4 -6 20 206
use INVX1  INVX1_190
timestamp 1651764895
transform -1 0 4744 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_217
timestamp 1651764895
transform 1 0 4744 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_91
timestamp 1651764895
transform -1 0 4840 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_77
timestamp 1651764895
transform 1 0 4840 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_84
timestamp 1651764895
transform -1 0 4936 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_139
timestamp 1651764895
transform 1 0 4936 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_204
timestamp 1651764895
transform 1 0 4968 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_191
timestamp 1651764895
transform -1 0 5080 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_207
timestamp 1651764895
transform 1 0 5080 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_26
timestamp 1651764895
transform 1 0 5144 0 -1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_195
timestamp 1651764895
transform -1 0 5304 0 -1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_104
timestamp 1651764895
transform 1 0 5304 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_218
timestamp 1651764895
transform 1 0 5368 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_219
timestamp 1651764895
transform -1 0 5496 0 -1 1810
box -4 -6 68 206
use AND2X2  AND2X2_57
timestamp 1651764895
transform 1 0 5496 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_191
timestamp 1651764895
transform 1 0 5560 0 -1 1810
box -4 -6 36 206
use INVX1  INVX1_192
timestamp 1651764895
transform 1 0 5592 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_205
timestamp 1651764895
transform 1 0 5624 0 -1 1810
box -4 -6 68 206
use NOR3X1  NOR3X1_22
timestamp 1651764895
transform 1 0 5688 0 -1 1810
box -4 -6 132 206
use XOR2X1  XOR2X1_16
timestamp 1651764895
transform -1 0 5928 0 -1 1810
box -4 -6 116 206
use DFFPOSX1  DFFPOSX1_11
timestamp 1651764895
transform 1 0 5928 0 -1 1810
box -4 -6 196 206
use BUFX2  BUFX2_28
timestamp 1651764895
transform 1 0 6120 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_309
timestamp 1651764895
transform 1 0 6168 0 -1 1810
box -4 -6 68 206
use FILL  FILL_9_1
timestamp 1651764895
transform -1 0 6248 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1651764895
transform -1 0 6264 0 -1 1810
box -4 -6 20 206
use AOI21X1  AOI21X1_39
timestamp 1651764895
transform 1 0 8 0 1 1810
box -4 -6 68 206
use AOI22X1  AOI22X1_6
timestamp 1651764895
transform 1 0 72 0 1 1810
box -4 -6 84 206
use AOI22X1  AOI22X1_11
timestamp 1651764895
transform 1 0 152 0 1 1810
box -4 -6 84 206
use INVX1  INVX1_127
timestamp 1651764895
transform 1 0 232 0 1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_71
timestamp 1651764895
transform 1 0 264 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_90
timestamp 1651764895
transform -1 0 376 0 1 1810
box -4 -6 52 206
use AND2X2  AND2X2_24
timestamp 1651764895
transform 1 0 376 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_118
timestamp 1651764895
transform 1 0 440 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_89
timestamp 1651764895
transform -1 0 536 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_25
timestamp 1651764895
transform 1 0 536 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_39
timestamp 1651764895
transform 1 0 584 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_65
timestamp 1651764895
transform 1 0 632 0 1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_5
timestamp 1651764895
transform 1 0 680 0 1 1810
box -4 -6 84 206
use NAND2X1  NAND2X1_38
timestamp 1651764895
transform 1 0 760 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_114
timestamp 1651764895
transform -1 0 856 0 1 1810
box -4 -6 52 206
use AND2X2  AND2X2_29
timestamp 1651764895
transform 1 0 856 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_28
timestamp 1651764895
transform -1 0 952 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_150
timestamp 1651764895
transform 1 0 952 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_149
timestamp 1651764895
transform 1 0 1016 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_134
timestamp 1651764895
transform -1 0 1144 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_85
timestamp 1651764895
transform 1 0 1144 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_131
timestamp 1651764895
transform 1 0 1208 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_176
timestamp 1651764895
transform 1 0 1272 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_135
timestamp 1651764895
transform -1 0 1400 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_150
timestamp 1651764895
transform 1 0 1400 0 1 1810
box -4 -6 36 206
use AOI22X1  AOI22X1_20
timestamp 1651764895
transform -1 0 1512 0 1 1810
box -4 -6 84 206
use AOI22X1  AOI22X1_19
timestamp 1651764895
transform -1 0 1592 0 1 1810
box -4 -6 84 206
use FILL  FILL_9_0_0
timestamp 1651764895
transform -1 0 1608 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1651764895
transform -1 0 1624 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1651764895
transform -1 0 1640 0 1 1810
box -4 -6 20 206
use NAND2X1  NAND2X1_146
timestamp 1651764895
transform -1 0 1688 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_147
timestamp 1651764895
transform 1 0 1688 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_136
timestamp 1651764895
transform 1 0 1736 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_94
timestamp 1651764895
transform 1 0 1800 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_182
timestamp 1651764895
transform 1 0 1864 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_194
timestamp 1651764895
transform -1 0 1960 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_193
timestamp 1651764895
transform 1 0 1960 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_189
timestamp 1651764895
transform -1 0 2088 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_97
timestamp 1651764895
transform 1 0 2088 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_191
timestamp 1651764895
transform -1 0 2216 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_96
timestamp 1651764895
transform 1 0 2216 0 1 1810
box -4 -6 68 206
use AND2X2  AND2X2_45
timestamp 1651764895
transform -1 0 2344 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_201
timestamp 1651764895
transform -1 0 2408 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_199
timestamp 1651764895
transform -1 0 2472 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_200
timestamp 1651764895
transform 1 0 2472 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_107
timestamp 1651764895
transform 1 0 2536 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_196
timestamp 1651764895
transform 1 0 2600 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_203
timestamp 1651764895
transform -1 0 2728 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_204
timestamp 1651764895
transform 1 0 2728 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_186
timestamp 1651764895
transform -1 0 2840 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_188
timestamp 1651764895
transform -1 0 2888 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_184
timestamp 1651764895
transform 1 0 2888 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_207
timestamp 1651764895
transform -1 0 3000 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_99
timestamp 1651764895
transform 1 0 3000 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_205
timestamp 1651764895
transform -1 0 3128 0 1 1810
box -4 -6 68 206
use FILL  FILL_9_1_0
timestamp 1651764895
transform 1 0 3128 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1651764895
transform 1 0 3144 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1651764895
transform 1 0 3160 0 1 1810
box -4 -6 20 206
use AOI21X1  AOI21X1_101
timestamp 1651764895
transform 1 0 3176 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_209
timestamp 1651764895
transform -1 0 3304 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_210
timestamp 1651764895
transform -1 0 3368 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_188
timestamp 1651764895
transform -1 0 3400 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_199
timestamp 1651764895
transform -1 0 3464 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_200
timestamp 1651764895
transform 1 0 3464 0 1 1810
box -4 -6 68 206
use OR2X2  OR2X2_18
timestamp 1651764895
transform 1 0 3528 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_170
timestamp 1651764895
transform -1 0 3656 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_131
timestamp 1651764895
transform 1 0 3656 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_130
timestamp 1651764895
transform 1 0 3720 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_103
timestamp 1651764895
transform 1 0 3784 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_54
timestamp 1651764895
transform 1 0 3832 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_211
timestamp 1651764895
transform -1 0 3944 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_102
timestamp 1651764895
transform 1 0 3944 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_190
timestamp 1651764895
transform -1 0 4056 0 1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_25
timestamp 1651764895
transform 1 0 4056 0 1 1810
box -4 -6 84 206
use OAI21X1  OAI21X1_201
timestamp 1651764895
transform 1 0 4136 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_202
timestamp 1651764895
transform 1 0 4200 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_189
timestamp 1651764895
transform -1 0 4296 0 1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_213
timestamp 1651764895
transform -1 0 4360 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_215
timestamp 1651764895
transform 1 0 4360 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_214
timestamp 1651764895
transform -1 0 4488 0 1 1810
box -4 -6 68 206
use AOI21X1  AOI21X1_103
timestamp 1651764895
transform 1 0 4488 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_159
timestamp 1651764895
transform -1 0 4600 0 1 1810
box -4 -6 52 206
use AOI22X1  AOI22X1_26
timestamp 1651764895
transform -1 0 4680 0 1 1810
box -4 -6 84 206
use FILL  FILL_9_2_0
timestamp 1651764895
transform 1 0 4680 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_1
timestamp 1651764895
transform 1 0 4696 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_2_2
timestamp 1651764895
transform 1 0 4712 0 1 1810
box -4 -6 20 206
use AND2X2  AND2X2_47
timestamp 1651764895
transform 1 0 4728 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_216
timestamp 1651764895
transform -1 0 4856 0 1 1810
box -4 -6 68 206
use AND2X2  AND2X2_56
timestamp 1651764895
transform 1 0 4856 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_89
timestamp 1651764895
transform -1 0 4984 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_82
timestamp 1651764895
transform 1 0 4984 0 1 1810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_20
timestamp 1651764895
transform -1 0 5144 0 1 1810
box -4 -6 116 206
use NAND2X1  NAND2X1_154
timestamp 1651764895
transform 1 0 5144 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_158
timestamp 1651764895
transform -1 0 5240 0 1 1810
box -4 -6 52 206
use OR2X2  OR2X2_17
timestamp 1651764895
transform -1 0 5304 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_208
timestamp 1651764895
transform 1 0 5304 0 1 1810
box -4 -6 68 206
use AOI22X1  AOI22X1_30
timestamp 1651764895
transform 1 0 5368 0 1 1810
box -4 -6 84 206
use NAND3X1  NAND3X1_273
timestamp 1651764895
transform -1 0 5512 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_223
timestamp 1651764895
transform -1 0 5544 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_251
timestamp 1651764895
transform -1 0 5608 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_252
timestamp 1651764895
transform 1 0 5608 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_276
timestamp 1651764895
transform -1 0 5736 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_277
timestamp 1651764895
transform -1 0 5800 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_136
timestamp 1651764895
transform 1 0 5800 0 1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_274
timestamp 1651764895
transform -1 0 5896 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_275
timestamp 1651764895
transform 1 0 5896 0 1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_278
timestamp 1651764895
transform 1 0 5960 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_250
timestamp 1651764895
transform -1 0 6072 0 1 1810
box -4 -6 52 206
use AOI21X1  AOI21X1_128
timestamp 1651764895
transform 1 0 6072 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_224
timestamp 1651764895
transform -1 0 6168 0 1 1810
box -4 -6 36 206
use AOI22X1  AOI22X1_37
timestamp 1651764895
transform 1 0 6168 0 1 1810
box -4 -6 84 206
use FILL  FILL_10_1
timestamp 1651764895
transform 1 0 6248 0 1 1810
box -4 -6 20 206
use NAND3X1  NAND3X1_73
timestamp 1651764895
transform -1 0 72 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_74
timestamp 1651764895
transform 1 0 72 0 -1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_78
timestamp 1651764895
transform -1 0 184 0 -1 2210
box -4 -6 52 206
use AND2X2  AND2X2_30
timestamp 1651764895
transform 1 0 184 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_64
timestamp 1651764895
transform 1 0 248 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_101
timestamp 1651764895
transform 1 0 312 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_145
timestamp 1651764895
transform 1 0 376 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_127
timestamp 1651764895
transform -1 0 504 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_148
timestamp 1651764895
transform -1 0 568 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_147
timestamp 1651764895
transform 1 0 568 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_129
timestamp 1651764895
transform 1 0 632 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_66
timestamp 1651764895
transform 1 0 696 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_128
timestamp 1651764895
transform 1 0 760 0 -1 2210
box -4 -6 68 206
use AOI22X1  AOI22X1_18
timestamp 1651764895
transform 1 0 824 0 -1 2210
box -4 -6 84 206
use INVX1  INVX1_181
timestamp 1651764895
transform 1 0 904 0 -1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_89
timestamp 1651764895
transform -1 0 1000 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_130
timestamp 1651764895
transform 1 0 1000 0 -1 2210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_21
timestamp 1651764895
transform 1 0 1064 0 -1 2210
box -4 -6 116 206
use NOR2X1  NOR2X1_87
timestamp 1651764895
transform -1 0 1224 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_75
timestamp 1651764895
transform 1 0 1224 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_74
timestamp 1651764895
transform 1 0 1272 0 -1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_120
timestamp 1651764895
transform -1 0 1384 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_139
timestamp 1651764895
transform -1 0 1448 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_140
timestamp 1651764895
transform 1 0 1448 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_118
timestamp 1651764895
transform 1 0 1512 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_0_0
timestamp 1651764895
transform 1 0 1576 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_1
timestamp 1651764895
transform 1 0 1592 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_0_2
timestamp 1651764895
transform 1 0 1608 0 -1 2210
box -4 -6 20 206
use NAND3X1  NAND3X1_133
timestamp 1651764895
transform 1 0 1624 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_121
timestamp 1651764895
transform -1 0 1752 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_151
timestamp 1651764895
transform 1 0 1752 0 -1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_132
timestamp 1651764895
transform 1 0 1784 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_119
timestamp 1651764895
transform 1 0 1848 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_169
timestamp 1651764895
transform 1 0 1912 0 -1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_93
timestamp 1651764895
transform -1 0 2024 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_186
timestamp 1651764895
transform 1 0 2024 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_92
timestamp 1651764895
transform -1 0 2152 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_187
timestamp 1651764895
transform 1 0 2152 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_188
timestamp 1651764895
transform -1 0 2280 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_190
timestamp 1651764895
transform 1 0 2280 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_109
timestamp 1651764895
transform 1 0 2344 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_220
timestamp 1651764895
transform -1 0 2472 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_171
timestamp 1651764895
transform -1 0 2520 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_183
timestamp 1651764895
transform 1 0 2520 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1651764895
transform 1 0 2568 0 -1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_278
timestamp 1651764895
transform 1 0 2600 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_279
timestamp 1651764895
transform -1 0 2696 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_181
timestamp 1651764895
transform 1 0 2696 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_219
timestamp 1651764895
transform -1 0 2808 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_185
timestamp 1651764895
transform 1 0 2808 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_168
timestamp 1651764895
transform 1 0 2856 0 -1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_202
timestamp 1651764895
transform 1 0 2904 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_182
timestamp 1651764895
transform -1 0 3016 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_107
timestamp 1651764895
transform -1 0 3064 0 -1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_206
timestamp 1651764895
transform 1 0 3064 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_1_0
timestamp 1651764895
transform -1 0 3144 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_1
timestamp 1651764895
transform -1 0 3160 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_1_2
timestamp 1651764895
transform -1 0 3176 0 -1 2210
box -4 -6 20 206
use NAND3X1  NAND3X1_208
timestamp 1651764895
transform -1 0 3240 0 -1 2210
box -4 -6 68 206
use AND2X2  AND2X2_48
timestamp 1651764895
transform 1 0 3240 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_217
timestamp 1651764895
transform 1 0 3304 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_124
timestamp 1651764895
transform -1 0 3384 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_172
timestamp 1651764895
transform -1 0 3448 0 -1 2210
box -4 -6 68 206
use AND2X2  AND2X2_40
timestamp 1651764895
transform 1 0 3448 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_36
timestamp 1651764895
transform -1 0 3544 0 -1 2210
box -4 -6 36 206
use INVX1  INVX1_43
timestamp 1651764895
transform -1 0 3576 0 -1 2210
box -4 -6 36 206
use OR2X2  OR2X2_20
timestamp 1651764895
transform 1 0 3576 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_171
timestamp 1651764895
transform -1 0 3704 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_163
timestamp 1651764895
transform -1 0 3752 0 -1 2210
box -4 -6 52 206
use NOR2X1  NOR2X1_94
timestamp 1651764895
transform 1 0 3752 0 -1 2210
box -4 -6 52 206
use AND2X2  AND2X2_41
timestamp 1651764895
transform 1 0 3800 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_172
timestamp 1651764895
transform 1 0 3864 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_174
timestamp 1651764895
transform 1 0 3896 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_213
timestamp 1651764895
transform 1 0 3960 0 -1 2210
box -4 -6 68 206
use AND2X2  AND2X2_46
timestamp 1651764895
transform 1 0 4024 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_212
timestamp 1651764895
transform -1 0 4152 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_264
timestamp 1651764895
transform -1 0 4216 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_125
timestamp 1651764895
transform -1 0 4280 0 -1 2210
box -4 -6 68 206
use AND2X2  AND2X2_53
timestamp 1651764895
transform 1 0 4280 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_207
timestamp 1651764895
transform 1 0 4344 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_247
timestamp 1651764895
transform 1 0 4392 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_248
timestamp 1651764895
transform 1 0 4456 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_268
timestamp 1651764895
transform 1 0 4520 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_266
timestamp 1651764895
transform 1 0 4584 0 -1 2210
box -4 -6 68 206
use FILL  FILL_10_2_0
timestamp 1651764895
transform -1 0 4664 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_1
timestamp 1651764895
transform -1 0 4680 0 -1 2210
box -4 -6 20 206
use FILL  FILL_10_2_2
timestamp 1651764895
transform -1 0 4696 0 -1 2210
box -4 -6 20 206
use NOR2X1  NOR2X1_67
timestamp 1651764895
transform -1 0 4744 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_115
timestamp 1651764895
transform 1 0 4744 0 -1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_126
timestamp 1651764895
transform -1 0 4840 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_196
timestamp 1651764895
transform 1 0 4840 0 -1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_88
timestamp 1651764895
transform -1 0 4952 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_267
timestamp 1651764895
transform -1 0 5016 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_126
timestamp 1651764895
transform 1 0 5016 0 -1 2210
box -4 -6 68 206
use AOI22X1  AOI22X1_29
timestamp 1651764895
transform 1 0 5080 0 -1 2210
box -4 -6 84 206
use INVX1  INVX1_254
timestamp 1651764895
transform 1 0 5160 0 -1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_156
timestamp 1651764895
transform -1 0 5256 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_269
timestamp 1651764895
transform -1 0 5320 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_249
timestamp 1651764895
transform 1 0 5320 0 -1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_250
timestamp 1651764895
transform 1 0 5384 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_272
timestamp 1651764895
transform -1 0 5512 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_270
timestamp 1651764895
transform 1 0 5512 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_255
timestamp 1651764895
transform 1 0 5576 0 -1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_127
timestamp 1651764895
transform -1 0 5688 0 -1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_271
timestamp 1651764895
transform -1 0 5752 0 -1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_157
timestamp 1651764895
transform 1 0 5752 0 -1 2210
box -4 -6 68 206
use INVX1  INVX1_255
timestamp 1651764895
transform -1 0 5848 0 -1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_251
timestamp 1651764895
transform 1 0 5848 0 -1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_305
timestamp 1651764895
transform 1 0 5896 0 -1 2210
box -4 -6 52 206
use INVX1  INVX1_257
timestamp 1651764895
transform 1 0 5944 0 -1 2210
box -4 -6 36 206
use AOI22X1  AOI22X1_38
timestamp 1651764895
transform 1 0 5976 0 -1 2210
box -4 -6 84 206
use NAND3X1  NAND3X1_333
timestamp 1651764895
transform 1 0 6056 0 -1 2210
box -4 -6 68 206
use AOI22X1  AOI22X1_39
timestamp 1651764895
transform 1 0 6120 0 -1 2210
box -4 -6 84 206
use AOI21X1  AOI21X1_159
timestamp 1651764895
transform 1 0 6200 0 -1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_116
timestamp 1651764895
transform -1 0 56 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_115
timestamp 1651764895
transform -1 0 104 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_117
timestamp 1651764895
transform -1 0 152 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_128
timestamp 1651764895
transform 1 0 152 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_102
timestamp 1651764895
transform -1 0 248 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_144
timestamp 1651764895
transform 1 0 248 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_125
timestamp 1651764895
transform -1 0 360 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_63
timestamp 1651764895
transform 1 0 360 0 1 2210
box -4 -6 68 206
use AOI22X1  AOI22X1_17
timestamp 1651764895
transform 1 0 424 0 1 2210
box -4 -6 84 206
use AND2X2  AND2X2_31
timestamp 1651764895
transform -1 0 568 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_86
timestamp 1651764895
transform 1 0 568 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_183
timestamp 1651764895
transform 1 0 632 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_144
timestamp 1651764895
transform 1 0 696 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_141
timestamp 1651764895
transform -1 0 808 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_143
timestamp 1651764895
transform 1 0 808 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_152
timestamp 1651764895
transform 1 0 872 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_139
timestamp 1651764895
transform 1 0 904 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_122
timestamp 1651764895
transform -1 0 1016 0 1 2210
box -4 -6 68 206
use AOI22X1  AOI22X1_23
timestamp 1651764895
transform 1 0 1016 0 1 2210
box -4 -6 84 206
use OAI21X1  OAI21X1_142
timestamp 1651764895
transform -1 0 1160 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_116
timestamp 1651764895
transform -1 0 1224 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_61
timestamp 1651764895
transform 1 0 1224 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_145
timestamp 1651764895
transform -1 0 1320 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_117
timestamp 1651764895
transform -1 0 1384 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_60
timestamp 1651764895
transform -1 0 1448 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_138
timestamp 1651764895
transform -1 0 1512 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_191
timestamp 1651764895
transform -1 0 1576 0 1 2210
box -4 -6 68 206
use FILL  FILL_11_0_0
timestamp 1651764895
transform 1 0 1576 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_1
timestamp 1651764895
transform 1 0 1592 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_0_2
timestamp 1651764895
transform 1 0 1608 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_192
timestamp 1651764895
transform 1 0 1624 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_185
timestamp 1651764895
transform -1 0 1752 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_110
timestamp 1651764895
transform 1 0 1752 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_182
timestamp 1651764895
transform 1 0 1816 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_222
timestamp 1651764895
transform 1 0 1880 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_175
timestamp 1651764895
transform -1 0 2008 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_175
timestamp 1651764895
transform -1 0 2056 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_180
timestamp 1651764895
transform -1 0 2104 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_213
timestamp 1651764895
transform 1 0 2104 0 1 2210
box -4 -6 36 206
use AOI21X1  AOI21X1_120
timestamp 1651764895
transform -1 0 2200 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_170
timestamp 1651764895
transform 1 0 2200 0 1 2210
box -4 -6 52 206
use OR2X2  OR2X2_21
timestamp 1651764895
transform 1 0 2248 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_245
timestamp 1651764895
transform -1 0 2376 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_251
timestamp 1651764895
transform -1 0 2440 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_246
timestamp 1651764895
transform -1 0 2504 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_201
timestamp 1651764895
transform 1 0 2504 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_252
timestamp 1651764895
transform 1 0 2536 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_249
timestamp 1651764895
transform 1 0 2600 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_250
timestamp 1651764895
transform -1 0 2728 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_254
timestamp 1651764895
transform -1 0 2792 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_216
timestamp 1651764895
transform -1 0 2824 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_253
timestamp 1651764895
transform 1 0 2824 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_255
timestamp 1651764895
transform 1 0 2888 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_187
timestamp 1651764895
transform 1 0 2952 0 1 2210
box -4 -6 52 206
use AOI21X1  AOI21X1_98
timestamp 1651764895
transform 1 0 3000 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_218
timestamp 1651764895
transform 1 0 3064 0 1 2210
box -4 -6 68 206
use FILL  FILL_11_1_0
timestamp 1651764895
transform 1 0 3128 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_1
timestamp 1651764895
transform 1 0 3144 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_1_2
timestamp 1651764895
transform 1 0 3160 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_171
timestamp 1651764895
transform 1 0 3176 0 1 2210
box -4 -6 68 206
use NOR2X1  NOR2X1_93
timestamp 1651764895
transform -1 0 3288 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_170
timestamp 1651764895
transform 1 0 3288 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_162
timestamp 1651764895
transform 1 0 3352 0 1 2210
box -4 -6 52 206
use OR2X2  OR2X2_19
timestamp 1651764895
transform -1 0 3464 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_214
timestamp 1651764895
transform -1 0 3528 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_127
timestamp 1651764895
transform -1 0 3576 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_210
timestamp 1651764895
transform -1 0 3624 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_215
timestamp 1651764895
transform 1 0 3624 0 1 2210
box -4 -6 52 206
use NAND2X1  NAND2X1_212
timestamp 1651764895
transform -1 0 3720 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_199
timestamp 1651764895
transform 1 0 3720 0 1 2210
box -4 -6 36 206
use NAND2X1  NAND2X1_214
timestamp 1651764895
transform 1 0 3752 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_225
timestamp 1651764895
transform -1 0 3864 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_200
timestamp 1651764895
transform -1 0 3896 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_224
timestamp 1651764895
transform 1 0 3896 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_213
timestamp 1651764895
transform 1 0 3960 0 1 2210
box -4 -6 52 206
use OAI21X1  OAI21X1_261
timestamp 1651764895
transform 1 0 4008 0 1 2210
box -4 -6 68 206
use AND2X2  AND2X2_61
timestamp 1651764895
transform 1 0 4072 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_249
timestamp 1651764895
transform 1 0 4136 0 1 2210
box -4 -6 52 206
use AND2X2  AND2X2_54
timestamp 1651764895
transform 1 0 4184 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_263
timestamp 1651764895
transform 1 0 4248 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_221
timestamp 1651764895
transform 1 0 4312 0 1 2210
box -4 -6 36 206
use AOI22X1  AOI22X1_28
timestamp 1651764895
transform 1 0 4344 0 1 2210
box -4 -6 84 206
use NOR2X1  NOR2X1_83
timestamp 1651764895
transform -1 0 4472 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_138
timestamp 1651764895
transform 1 0 4472 0 1 2210
box -4 -6 36 206
use NOR2X1  NOR2X1_68
timestamp 1651764895
transform -1 0 4552 0 1 2210
box -4 -6 52 206
use INVX1  INVX1_116
timestamp 1651764895
transform 1 0 4552 0 1 2210
box -4 -6 36 206
use OAI21X1  OAI21X1_166
timestamp 1651764895
transform 1 0 4584 0 1 2210
box -4 -6 68 206
use FILL  FILL_11_2_0
timestamp 1651764895
transform 1 0 4648 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_1
timestamp 1651764895
transform 1 0 4664 0 1 2210
box -4 -6 20 206
use FILL  FILL_11_2_2
timestamp 1651764895
transform 1 0 4680 0 1 2210
box -4 -6 20 206
use OAI21X1  OAI21X1_127
timestamp 1651764895
transform 1 0 4696 0 1 2210
box -4 -6 68 206
use OAI22X1  OAI22X1_5
timestamp 1651764895
transform 1 0 4760 0 1 2210
box -4 -6 84 206
use XOR2X1  XOR2X1_9
timestamp 1651764895
transform -1 0 4952 0 1 2210
box -4 -6 116 206
use AND2X2  AND2X2_55
timestamp 1651764895
transform -1 0 5016 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_206
timestamp 1651764895
transform 1 0 5016 0 1 2210
box -4 -6 52 206
use OR2X2  OR2X2_25
timestamp 1651764895
transform -1 0 5128 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_205
timestamp 1651764895
transform 1 0 5128 0 1 2210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_31
timestamp 1651764895
transform 1 0 5176 0 1 2210
box -4 -6 116 206
use NAND2X1  NAND2X1_252
timestamp 1651764895
transform 1 0 5288 0 1 2210
box -4 -6 52 206
use AND2X2  AND2X2_59
timestamp 1651764895
transform 1 0 5336 0 1 2210
box -4 -6 68 206
use AND2X2  AND2X2_58
timestamp 1651764895
transform -1 0 5464 0 1 2210
box -4 -6 68 206
use NAND2X1  NAND2X1_204
timestamp 1651764895
transform -1 0 5512 0 1 2210
box -4 -6 52 206
use NAND3X1  NAND3X1_331
timestamp 1651764895
transform -1 0 5576 0 1 2210
box -4 -6 68 206
use AOI21X1  AOI21X1_158
timestamp 1651764895
transform 1 0 5576 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_307
timestamp 1651764895
transform 1 0 5640 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_306
timestamp 1651764895
transform 1 0 5704 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_334
timestamp 1651764895
transform 1 0 5768 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_332
timestamp 1651764895
transform -1 0 5896 0 1 2210
box -4 -6 68 206
use NAND3X1  NAND3X1_335
timestamp 1651764895
transform -1 0 5960 0 1 2210
box -4 -6 68 206
use INVX1  INVX1_256
timestamp 1651764895
transform -1 0 5992 0 1 2210
box -4 -6 36 206
use NAND3X1  NAND3X1_336
timestamp 1651764895
transform 1 0 5992 0 1 2210
box -4 -6 68 206
use OAI21X1  OAI21X1_366
timestamp 1651764895
transform 1 0 6056 0 1 2210
box -4 -6 68 206
use XNOR2X1  XNOR2X1_37
timestamp 1651764895
transform 1 0 6120 0 1 2210
box -4 -6 116 206
use FILL  FILL_12_1
timestamp 1651764895
transform 1 0 6232 0 1 2210
box -4 -6 20 206
use FILL  FILL_12_2
timestamp 1651764895
transform 1 0 6248 0 1 2210
box -4 -6 20 206
use BUFX2  BUFX2_17
timestamp 1651764895
transform 1 0 8 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_14
timestamp 1651764895
transform 1 0 56 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_124
timestamp 1651764895
transform 1 0 104 0 -1 2610
box -4 -6 68 206
use BUFX2  BUFX2_16
timestamp 1651764895
transform 1 0 168 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_15
timestamp 1651764895
transform 1 0 216 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_123
timestamp 1651764895
transform -1 0 328 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_154
timestamp 1651764895
transform -1 0 360 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_186
timestamp 1651764895
transform 1 0 360 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_126
timestamp 1651764895
transform -1 0 488 0 -1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_24
timestamp 1651764895
transform -1 0 568 0 -1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_146
timestamp 1651764895
transform -1 0 632 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_15
timestamp 1651764895
transform 1 0 632 0 -1 2610
box -4 -6 36 206
use AND2X2  AND2X2_38
timestamp 1651764895
transform 1 0 664 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_180
timestamp 1651764895
transform -1 0 792 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_178
timestamp 1651764895
transform -1 0 856 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_112
timestamp 1651764895
transform 1 0 856 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_189
timestamp 1651764895
transform -1 0 984 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_190
timestamp 1651764895
transform 1 0 984 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_138
timestamp 1651764895
transform 1 0 1048 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_176
timestamp 1651764895
transform -1 0 1144 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_180
timestamp 1651764895
transform 1 0 1144 0 -1 2610
box -4 -6 36 206
use XNOR2X1  XNOR2X1_28
timestamp 1651764895
transform -1 0 1288 0 -1 2610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_27
timestamp 1651764895
transform -1 0 1400 0 -1 2610
box -4 -6 116 206
use NAND3X1  NAND3X1_179
timestamp 1651764895
transform -1 0 1464 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_91
timestamp 1651764895
transform 1 0 1464 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_227
timestamp 1651764895
transform 1 0 1528 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_0_0
timestamp 1651764895
transform 1 0 1592 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_1
timestamp 1651764895
transform 1 0 1608 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_0_2
timestamp 1651764895
transform 1 0 1624 0 -1 2610
box -4 -6 20 206
use OAI21X1  OAI21X1_137
timestamp 1651764895
transform 1 0 1640 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_137
timestamp 1651764895
transform -1 0 1752 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_149
timestamp 1651764895
transform -1 0 1784 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_147
timestamp 1651764895
transform -1 0 1816 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_177
timestamp 1651764895
transform 1 0 1816 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_181
timestamp 1651764895
transform 1 0 1880 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_90
timestamp 1651764895
transform -1 0 2008 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_115
timestamp 1651764895
transform 1 0 2008 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_212
timestamp 1651764895
transform 1 0 2072 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_182
timestamp 1651764895
transform 1 0 2104 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_184
timestamp 1651764895
transform -1 0 2232 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_174
timestamp 1651764895
transform 1 0 2232 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_181
timestamp 1651764895
transform 1 0 2296 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_176
timestamp 1651764895
transform 1 0 2360 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_172
timestamp 1651764895
transform 1 0 2392 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_175
timestamp 1651764895
transform 1 0 2456 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_173
timestamp 1651764895
transform 1 0 2488 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_183
timestamp 1651764895
transform 1 0 2552 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_221
timestamp 1651764895
transform -1 0 2664 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_240
timestamp 1651764895
transform -1 0 2728 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_239
timestamp 1651764895
transform 1 0 2728 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_215
timestamp 1651764895
transform 1 0 2792 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_244
timestamp 1651764895
transform 1 0 2824 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_248
timestamp 1651764895
transform -1 0 2952 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_243
timestamp 1651764895
transform 1 0 2952 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_151
timestamp 1651764895
transform -1 0 3080 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_1_0
timestamp 1651764895
transform 1 0 3080 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_1
timestamp 1651764895
transform 1 0 3096 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_1_2
timestamp 1651764895
transform 1 0 3112 0 -1 2610
box -4 -6 20 206
use NAND3X1  NAND3X1_247
timestamp 1651764895
transform 1 0 3128 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_108
timestamp 1651764895
transform -1 0 3256 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_280
timestamp 1651764895
transform 1 0 3256 0 -1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_32
timestamp 1651764895
transform -1 0 3384 0 -1 2610
box -4 -6 84 206
use NAND2X1  NAND2X1_239
timestamp 1651764895
transform -1 0 3432 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_241
timestamp 1651764895
transform 1 0 3432 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_241
timestamp 1651764895
transform 1 0 3480 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_242
timestamp 1651764895
transform -1 0 3592 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_123
timestamp 1651764895
transform 1 0 3592 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_211
timestamp 1651764895
transform 1 0 3656 0 -1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_243
timestamp 1651764895
transform -1 0 3768 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_217
timestamp 1651764895
transform 1 0 3768 0 -1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_244
timestamp 1651764895
transform 1 0 3800 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_260
timestamp 1651764895
transform -1 0 3912 0 -1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_31
timestamp 1651764895
transform -1 0 3992 0 -1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_217
timestamp 1651764895
transform 1 0 3992 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_65
timestamp 1651764895
transform -1 0 4088 0 -1 2610
box -4 -6 36 206
use INVX1  INVX1_198
timestamp 1651764895
transform 1 0 4088 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_223
timestamp 1651764895
transform 1 0 4120 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_22
timestamp 1651764895
transform -1 0 4216 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_261
timestamp 1651764895
transform -1 0 4280 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_247
timestamp 1651764895
transform 1 0 4280 0 -1 2610
box -4 -6 52 206
use AOI21X1  AOI21X1_124
timestamp 1651764895
transform 1 0 4328 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_220
timestamp 1651764895
transform 1 0 4392 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_265
timestamp 1651764895
transform -1 0 4488 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_248
timestamp 1651764895
transform -1 0 4536 0 -1 2610
box -4 -6 52 206
use AND2X2  AND2X2_65
timestamp 1651764895
transform -1 0 4600 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_245
timestamp 1651764895
transform -1 0 4664 0 -1 2610
box -4 -6 68 206
use FILL  FILL_12_2_0
timestamp 1651764895
transform 1 0 4664 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_1
timestamp 1651764895
transform 1 0 4680 0 -1 2610
box -4 -6 20 206
use FILL  FILL_12_2_2
timestamp 1651764895
transform 1 0 4696 0 -1 2610
box -4 -6 20 206
use OAI21X1  OAI21X1_246
timestamp 1651764895
transform 1 0 4712 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_222
timestamp 1651764895
transform -1 0 4808 0 -1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_262
timestamp 1651764895
transform 1 0 4808 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_266
timestamp 1651764895
transform -1 0 4920 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_265
timestamp 1651764895
transform 1 0 4920 0 -1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_155
timestamp 1651764895
transform 1 0 4984 0 -1 2610
box -4 -6 68 206
use INVX1  INVX1_253
timestamp 1651764895
transform 1 0 5048 0 -1 2610
box -4 -6 36 206
use NOR2X1  NOR2X1_90
timestamp 1651764895
transform 1 0 5080 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_168
timestamp 1651764895
transform 1 0 5128 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_167
timestamp 1651764895
transform -1 0 5224 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_211
timestamp 1651764895
transform 1 0 5224 0 -1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_92
timestamp 1651764895
transform 1 0 5288 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_170
timestamp 1651764895
transform 1 0 5336 0 -1 2610
box -4 -6 36 206
use OAI21X1  OAI21X1_168
timestamp 1651764895
transform 1 0 5368 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_157
timestamp 1651764895
transform 1 0 5432 0 -1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_221
timestamp 1651764895
transform -1 0 5544 0 -1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_264
timestamp 1651764895
transform -1 0 5592 0 -1 2610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_24
timestamp 1651764895
transform -1 0 5704 0 -1 2610
box -4 -6 116 206
use NAND2X1  NAND2X1_262
timestamp 1651764895
transform 1 0 5704 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_263
timestamp 1651764895
transform -1 0 5800 0 -1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_261
timestamp 1651764895
transform -1 0 5848 0 -1 2610
box -4 -6 52 206
use INVX1  INVX1_233
timestamp 1651764895
transform 1 0 5848 0 -1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_198
timestamp 1651764895
transform 1 0 5880 0 -1 2610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_25
timestamp 1651764895
transform 1 0 5928 0 -1 2610
box -4 -6 116 206
use OAI21X1  OAI21X1_305
timestamp 1651764895
transform -1 0 6104 0 -1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_304
timestamp 1651764895
transform 1 0 6104 0 -1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_330
timestamp 1651764895
transform 1 0 6168 0 -1 2610
box -4 -6 68 206
use FILL  FILL_13_1
timestamp 1651764895
transform -1 0 6248 0 -1 2610
box -4 -6 20 206
use FILL  FILL_13_2
timestamp 1651764895
transform -1 0 6264 0 -1 2610
box -4 -6 20 206
use BUFX2  BUFX2_4
timestamp 1651764895
transform 1 0 8 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1651764895
transform 1 0 56 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_145
timestamp 1651764895
transform -1 0 152 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_3
timestamp 1651764895
transform 1 0 152 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_2
timestamp 1651764895
transform 1 0 200 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_143
timestamp 1651764895
transform 1 0 248 0 1 2610
box -4 -6 52 206
use AND2X2  AND2X2_37
timestamp 1651764895
transform 1 0 296 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_97
timestamp 1651764895
transform 1 0 360 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_142
timestamp 1651764895
transform 1 0 408 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_10
timestamp 1651764895
transform 1 0 456 0 1 2610
box -4 -6 36 206
use AND2X2  AND2X2_43
timestamp 1651764895
transform 1 0 488 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_188
timestamp 1651764895
transform 1 0 552 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_179
timestamp 1651764895
transform 1 0 616 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_187
timestamp 1651764895
transform 1 0 664 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_176
timestamp 1651764895
transform -1 0 792 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_88
timestamp 1651764895
transform 1 0 792 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_178
timestamp 1651764895
transform -1 0 904 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_178
timestamp 1651764895
transform 1 0 904 0 1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_87
timestamp 1651764895
transform 1 0 936 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_84
timestamp 1651764895
transform -1 0 1048 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_140
timestamp 1651764895
transform 1 0 1048 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_185
timestamp 1651764895
transform -1 0 1160 0 1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_10
timestamp 1651764895
transform 1 0 1160 0 1 2610
box -4 -6 84 206
use OAI22X1  OAI22X1_7
timestamp 1651764895
transform 1 0 1240 0 1 2610
box -4 -6 84 206
use NOR2X1  NOR2X1_86
timestamp 1651764895
transform -1 0 1368 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_108
timestamp 1651764895
transform 1 0 1368 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_136
timestamp 1651764895
transform 1 0 1416 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_136
timestamp 1651764895
transform 1 0 1480 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_179
timestamp 1651764895
transform -1 0 1592 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_0_0
timestamp 1651764895
transform -1 0 1608 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_1
timestamp 1651764895
transform -1 0 1624 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_0_2
timestamp 1651764895
transform -1 0 1640 0 1 2610
box -4 -6 20 206
use NAND2X1  NAND2X1_174
timestamp 1651764895
transform -1 0 1688 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_180
timestamp 1651764895
transform 1 0 1688 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_205
timestamp 1651764895
transform 1 0 1752 0 1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_111
timestamp 1651764895
transform 1 0 1784 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_96
timestamp 1651764895
transform -1 0 1896 0 1 2610
box -4 -6 52 206
use OR2X2  OR2X2_22
timestamp 1651764895
transform 1 0 1896 0 1 2610
box -4 -6 68 206
use AND2X2  AND2X2_42
timestamp 1651764895
transform 1 0 1960 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_95
timestamp 1651764895
transform -1 0 2072 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_240
timestamp 1651764895
transform -1 0 2136 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_131
timestamp 1651764895
transform -1 0 2200 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_238
timestamp 1651764895
transform 1 0 2200 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_239
timestamp 1651764895
transform -1 0 2328 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_122
timestamp 1651764895
transform 1 0 2328 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_242
timestamp 1651764895
transform -1 0 2456 0 1 2610
box -4 -6 68 206
use AOI21X1  AOI21X1_130
timestamp 1651764895
transform 1 0 2456 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_266
timestamp 1651764895
transform 1 0 2520 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_202
timestamp 1651764895
transform 1 0 2584 0 1 2610
box -4 -6 36 206
use INVX1  INVX1_248
timestamp 1651764895
transform 1 0 2616 0 1 2610
box -4 -6 36 206
use AOI21X1  AOI21X1_150
timestamp 1651764895
transform -1 0 2712 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_242
timestamp 1651764895
transform -1 0 2776 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_243
timestamp 1651764895
transform 1 0 2776 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_354
timestamp 1651764895
transform 1 0 2824 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_257
timestamp 1651764895
transform -1 0 2952 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_258
timestamp 1651764895
transform -1 0 3016 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_218
timestamp 1651764895
transform 1 0 3016 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_259
timestamp 1651764895
transform -1 0 3128 0 1 2610
box -4 -6 68 206
use FILL  FILL_13_1_0
timestamp 1651764895
transform 1 0 3128 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_1
timestamp 1651764895
transform 1 0 3144 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_1_2
timestamp 1651764895
transform 1 0 3160 0 1 2610
box -4 -6 20 206
use NAND3X1  NAND3X1_256
timestamp 1651764895
transform 1 0 3176 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_240
timestamp 1651764895
transform -1 0 3288 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_161
timestamp 1651764895
transform -1 0 3336 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_215
timestamp 1651764895
transform 1 0 3336 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_216
timestamp 1651764895
transform -1 0 3464 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_262
timestamp 1651764895
transform 1 0 3464 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_273
timestamp 1651764895
transform 1 0 3528 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_236
timestamp 1651764895
transform -1 0 3608 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_271
timestamp 1651764895
transform 1 0 3608 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_237
timestamp 1651764895
transform 1 0 3656 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_274
timestamp 1651764895
transform -1 0 3736 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_272
timestamp 1651764895
transform 1 0 3736 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_283
timestamp 1651764895
transform -1 0 3848 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_317
timestamp 1651764895
transform -1 0 3912 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_238
timestamp 1651764895
transform 1 0 3912 0 1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_318
timestamp 1651764895
transform 1 0 3944 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_284
timestamp 1651764895
transform 1 0 4008 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_301
timestamp 1651764895
transform 1 0 4072 0 1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_33
timestamp 1651764895
transform 1 0 4120 0 1 2610
box -4 -6 84 206
use NAND3X1  NAND3X1_320
timestamp 1651764895
transform -1 0 4264 0 1 2610
box -4 -6 68 206
use AOI22X1  AOI22X1_34
timestamp 1651764895
transform -1 0 4344 0 1 2610
box -4 -6 84 206
use OAI21X1  OAI21X1_302
timestamp 1651764895
transform 1 0 4344 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_303
timestamp 1651764895
transform 1 0 4408 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_322
timestamp 1651764895
transform -1 0 4536 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_326
timestamp 1651764895
transform 1 0 4536 0 1 2610
box -4 -6 68 206
use NOR2X1  NOR2X1_91
timestamp 1651764895
transform -1 0 4648 0 1 2610
box -4 -6 52 206
use FILL  FILL_13_2_0
timestamp 1651764895
transform 1 0 4648 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_1
timestamp 1651764895
transform 1 0 4664 0 1 2610
box -4 -6 20 206
use FILL  FILL_13_2_2
timestamp 1651764895
transform 1 0 4680 0 1 2610
box -4 -6 20 206
use INVX1  INVX1_169
timestamp 1651764895
transform 1 0 4696 0 1 2610
box -4 -6 36 206
use INVX1  INVX1_167
timestamp 1651764895
transform -1 0 4760 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_124
timestamp 1651764895
transform 1 0 4760 0 1 2610
box -4 -6 52 206
use OAI21X1  OAI21X1_212
timestamp 1651764895
transform 1 0 4808 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_200
timestamp 1651764895
transform -1 0 4920 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_201
timestamp 1651764895
transform 1 0 4920 0 1 2610
box -4 -6 52 206
use OR2X2  OR2X2_23
timestamp 1651764895
transform 1 0 4968 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_202
timestamp 1651764895
transform 1 0 5032 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_196
timestamp 1651764895
transform -1 0 5112 0 1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_325
timestamp 1651764895
transform -1 0 5176 0 1 2610
box -4 -6 68 206
use NAND3X1  NAND3X1_282
timestamp 1651764895
transform -1 0 5240 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_234
timestamp 1651764895
transform 1 0 5240 0 1 2610
box -4 -6 36 206
use NAND3X1  NAND3X1_324
timestamp 1651764895
transform 1 0 5272 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_303
timestamp 1651764895
transform 1 0 5336 0 1 2610
box -4 -6 52 206
use AOI22X1  AOI22X1_36
timestamp 1651764895
transform 1 0 5384 0 1 2610
box -4 -6 84 206
use NAND3X1  NAND3X1_323
timestamp 1651764895
transform 1 0 5464 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_254
timestamp 1651764895
transform -1 0 5592 0 1 2610
box -4 -6 68 206
use OR2X2  OR2X2_24
timestamp 1651764895
transform -1 0 5656 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_203
timestamp 1651764895
transform -1 0 5704 0 1 2610
box -4 -6 52 206
use NAND3X1  NAND3X1_281
timestamp 1651764895
transform 1 0 5704 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_210
timestamp 1651764895
transform -1 0 5832 0 1 2610
box -4 -6 68 206
use INVX1  INVX1_193
timestamp 1651764895
transform 1 0 5832 0 1 2610
box -4 -6 36 206
use NAND2X1  NAND2X1_253
timestamp 1651764895
transform 1 0 5864 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_195
timestamp 1651764895
transform 1 0 5912 0 1 2610
box -4 -6 36 206
use OR2X2  OR2X2_27
timestamp 1651764895
transform 1 0 5944 0 1 2610
box -4 -6 68 206
use OAI21X1  OAI21X1_253
timestamp 1651764895
transform -1 0 6072 0 1 2610
box -4 -6 68 206
use NAND2X1  NAND2X1_155
timestamp 1651764895
transform -1 0 6120 0 1 2610
box -4 -6 52 206
use NAND2X1  NAND2X1_254
timestamp 1651764895
transform -1 0 6168 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_29
timestamp 1651764895
transform 1 0 6168 0 1 2610
box -4 -6 52 206
use INVX1  INVX1_225
timestamp 1651764895
transform -1 0 6248 0 1 2610
box -4 -6 36 206
use FILL  FILL_14_1
timestamp 1651764895
transform 1 0 6248 0 1 2610
box -4 -6 20 206
use NAND2X1  NAND2X1_512
timestamp 1651764895
transform -1 0 56 0 -1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_70
timestamp 1651764895
transform -1 0 168 0 -1 3010
box -4 -6 116 206
use NAND2X1  NAND2X1_468
timestamp 1651764895
transform -1 0 216 0 -1 3010
box -4 -6 52 206
use AOI22X1  AOI22X1_40
timestamp 1651764895
transform 1 0 216 0 -1 3010
box -4 -6 84 206
use AND2X2  AND2X2_76
timestamp 1651764895
transform 1 0 296 0 -1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_147
timestamp 1651764895
transform -1 0 408 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_292
timestamp 1651764895
transform -1 0 456 0 -1 3010
box -4 -6 52 206
use AND2X2  AND2X2_44
timestamp 1651764895
transform 1 0 456 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_71
timestamp 1651764895
transform -1 0 552 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_233
timestamp 1651764895
transform -1 0 600 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_291
timestamp 1651764895
transform -1 0 648 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_208
timestamp 1651764895
transform 1 0 648 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_234
timestamp 1651764895
transform 1 0 680 0 -1 3010
box -4 -6 52 206
use OAI22X1  OAI22X1_6
timestamp 1651764895
transform 1 0 728 0 -1 3010
box -4 -6 84 206
use AOI22X1  AOI22X1_27
timestamp 1651764895
transform 1 0 808 0 -1 3010
box -4 -6 84 206
use NAND3X1  NAND3X1_177
timestamp 1651764895
transform 1 0 888 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_148
timestamp 1651764895
transform -1 0 984 0 -1 3010
box -4 -6 36 206
use INVX1  INVX1_46
timestamp 1651764895
transform 1 0 984 0 -1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_184
timestamp 1651764895
transform 1 0 1016 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_144
timestamp 1651764895
transform 1 0 1080 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_177
timestamp 1651764895
transform 1 0 1112 0 -1 3010
box -4 -6 52 206
use XOR2X1  XOR2X1_14
timestamp 1651764895
transform 1 0 1160 0 -1 3010
box -4 -6 116 206
use XNOR2X1  XNOR2X1_32
timestamp 1651764895
transform -1 0 1384 0 -1 3010
box -4 -6 116 206
use OAI21X1  OAI21X1_178
timestamp 1651764895
transform -1 0 1448 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_232
timestamp 1651764895
transform -1 0 1512 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_236
timestamp 1651764895
transform 1 0 1512 0 -1 3010
box -4 -6 68 206
use FILL  FILL_14_0_0
timestamp 1651764895
transform 1 0 1576 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_1
timestamp 1651764895
transform 1 0 1592 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_0_2
timestamp 1651764895
transform 1 0 1608 0 -1 3010
box -4 -6 20 206
use OAI21X1  OAI21X1_235
timestamp 1651764895
transform 1 0 1624 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_235
timestamp 1651764895
transform -1 0 1752 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_231
timestamp 1651764895
transform -1 0 1816 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_132
timestamp 1651764895
transform -1 0 1880 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_119
timestamp 1651764895
transform 1 0 1880 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_236
timestamp 1651764895
transform 1 0 1944 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_118
timestamp 1651764895
transform 1 0 2008 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_237
timestamp 1651764895
transform -1 0 2136 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_237
timestamp 1651764895
transform -1 0 2200 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_238
timestamp 1651764895
transform 1 0 2200 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_267
timestamp 1651764895
transform -1 0 2328 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_121
timestamp 1651764895
transform 1 0 2328 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_241
timestamp 1651764895
transform 1 0 2392 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_214
timestamp 1651764895
transform -1 0 2488 0 -1 3010
box -4 -6 36 206
use INVX1  INVX1_247
timestamp 1651764895
transform 1 0 2488 0 -1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_145
timestamp 1651764895
transform 1 0 2520 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_294
timestamp 1651764895
transform -1 0 2648 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_295
timestamp 1651764895
transform 1 0 2648 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_304
timestamp 1651764895
transform 1 0 2712 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_305
timestamp 1651764895
transform -1 0 2840 0 -1 3010
box -4 -6 68 206
use AOI22X1  AOI22X1_41
timestamp 1651764895
transform 1 0 2840 0 -1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_347
timestamp 1651764895
transform -1 0 2968 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_307
timestamp 1651764895
transform -1 0 3032 0 -1 3010
box -4 -6 68 206
use AND2X2  AND2X2_78
timestamp 1651764895
transform -1 0 3096 0 -1 3010
box -4 -6 68 206
use FILL  FILL_14_1_0
timestamp 1651764895
transform -1 0 3112 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_1
timestamp 1651764895
transform -1 0 3128 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_1_2
timestamp 1651764895
transform -1 0 3144 0 -1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_296
timestamp 1651764895
transform -1 0 3192 0 -1 3010
box -4 -6 52 206
use AND2X2  AND2X2_64
timestamp 1651764895
transform 1 0 3192 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_245
timestamp 1651764895
transform -1 0 3304 0 -1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_117
timestamp 1651764895
transform 1 0 3304 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_208
timestamp 1651764895
transform 1 0 3352 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_235
timestamp 1651764895
transform 1 0 3400 0 -1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_277
timestamp 1651764895
transform 1 0 3432 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_269
timestamp 1651764895
transform 1 0 3480 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_209
timestamp 1651764895
transform -1 0 3576 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_263
timestamp 1651764895
transform 1 0 3576 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_268
timestamp 1651764895
transform 1 0 3640 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_267
timestamp 1651764895
transform 1 0 3688 0 -1 3010
box -4 -6 52 206
use OR2X2  OR2X2_31
timestamp 1651764895
transform 1 0 3736 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_320
timestamp 1651764895
transform -1 0 3864 0 -1 3010
box -4 -6 68 206
use OR2X2  OR2X2_28
timestamp 1651764895
transform 1 0 3864 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_270
timestamp 1651764895
transform -1 0 3976 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_264
timestamp 1651764895
transform -1 0 4040 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_319
timestamp 1651764895
transform 1 0 4040 0 -1 3010
box -4 -6 68 206
use AND2X2  AND2X2_72
timestamp 1651764895
transform 1 0 4104 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_316
timestamp 1651764895
transform -1 0 4232 0 -1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_319
timestamp 1651764895
transform 1 0 4232 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_301
timestamp 1651764895
transform -1 0 4360 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_300
timestamp 1651764895
transform 1 0 4360 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_302
timestamp 1651764895
transform 1 0 4424 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_321
timestamp 1651764895
transform 1 0 4472 0 -1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_161
timestamp 1651764895
transform 1 0 4536 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_270
timestamp 1651764895
transform -1 0 4632 0 -1 3010
box -4 -6 36 206
use FILL  FILL_14_2_0
timestamp 1651764895
transform 1 0 4632 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_1
timestamp 1651764895
transform 1 0 4648 0 -1 3010
box -4 -6 20 206
use FILL  FILL_14_2_2
timestamp 1651764895
transform 1 0 4664 0 -1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_311
timestamp 1651764895
transform 1 0 4680 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_534
timestamp 1651764895
transform -1 0 4776 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_536
timestamp 1651764895
transform -1 0 4824 0 -1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_79
timestamp 1651764895
transform -1 0 4936 0 -1 3010
box -4 -6 116 206
use INVX1  INVX1_114
timestamp 1651764895
transform -1 0 4968 0 -1 3010
box -4 -6 36 206
use INVX1  INVX1_197
timestamp 1651764895
transform -1 0 5000 0 -1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_222
timestamp 1651764895
transform -1 0 5064 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_257
timestamp 1651764895
transform -1 0 5112 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_258
timestamp 1651764895
transform -1 0 5176 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_229
timestamp 1651764895
transform -1 0 5208 0 -1 3010
box -4 -6 36 206
use NOR2X1  NOR2X1_101
timestamp 1651764895
transform 1 0 5208 0 -1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_30
timestamp 1651764895
transform 1 0 5256 0 -1 3010
box -4 -6 116 206
use NAND2X1  NAND2X1_156
timestamp 1651764895
transform 1 0 5368 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_436
timestamp 1651764895
transform -1 0 5464 0 -1 3010
box -4 -6 52 206
use INVX1  INVX1_295
timestamp 1651764895
transform 1 0 5464 0 -1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_190
timestamp 1651764895
transform -1 0 5560 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_265
timestamp 1651764895
transform -1 0 5608 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_310
timestamp 1651764895
transform 1 0 5608 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_327
timestamp 1651764895
transform 1 0 5656 0 -1 3010
box -4 -6 68 206
use AOI22X1  AOI22X1_35
timestamp 1651764895
transform -1 0 5800 0 -1 3010
box -4 -6 84 206
use AND2X2  AND2X2_67
timestamp 1651764895
transform -1 0 5864 0 -1 3010
box -4 -6 68 206
use INVX1  INVX1_194
timestamp 1651764895
transform 1 0 5864 0 -1 3010
box -4 -6 36 206
use NOR2X1  NOR2X1_100
timestamp 1651764895
transform -1 0 5944 0 -1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_209
timestamp 1651764895
transform 1 0 5944 0 -1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_255
timestamp 1651764895
transform -1 0 6072 0 -1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_256
timestamp 1651764895
transform -1 0 6120 0 -1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_199
timestamp 1651764895
transform -1 0 6168 0 -1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_329
timestamp 1651764895
transform 1 0 6168 0 -1 3010
box -4 -6 68 206
use FILL  FILL_15_1
timestamp 1651764895
transform -1 0 6248 0 -1 3010
box -4 -6 20 206
use FILL  FILL_15_2
timestamp 1651764895
transform -1 0 6264 0 -1 3010
box -4 -6 20 206
use XNOR2X1  XNOR2X1_71
timestamp 1651764895
transform 1 0 8 0 1 3010
box -4 -6 116 206
use NAND2X1  NAND2X1_511
timestamp 1651764895
transform -1 0 168 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_470
timestamp 1651764895
transform -1 0 216 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_469
timestamp 1651764895
transform -1 0 264 0 1 3010
box -4 -6 52 206
use AND2X2  AND2X2_63
timestamp 1651764895
transform 1 0 264 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_235
timestamp 1651764895
transform 1 0 328 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_125
timestamp 1651764895
transform -1 0 424 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_105
timestamp 1651764895
transform -1 0 472 0 1 3010
box -4 -6 52 206
use AND2X2  AND2X2_51
timestamp 1651764895
transform 1 0 472 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_231
timestamp 1651764895
transform 1 0 536 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_153
timestamp 1651764895
transform -1 0 632 0 1 3010
box -4 -6 36 206
use NOR3X1  NOR3X1_21
timestamp 1651764895
transform -1 0 760 0 1 3010
box -4 -6 132 206
use NAND2X1  NAND2X1_236
timestamp 1651764895
transform 1 0 760 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_230
timestamp 1651764895
transform 1 0 808 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_279
timestamp 1651764895
transform 1 0 872 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_209
timestamp 1651764895
transform 1 0 936 0 1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_134
timestamp 1651764895
transform -1 0 1032 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_114
timestamp 1651764895
transform 1 0 1032 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_228
timestamp 1651764895
transform 1 0 1096 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_233
timestamp 1651764895
transform 1 0 1160 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_234
timestamp 1651764895
transform 1 0 1224 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_232
timestamp 1651764895
transform -1 0 1352 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_117
timestamp 1651764895
transform 1 0 1352 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_211
timestamp 1651764895
transform 1 0 1416 0 1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_113
timestamp 1651764895
transform 1 0 1448 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_229
timestamp 1651764895
transform -1 0 1576 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_0_0
timestamp 1651764895
transform 1 0 1576 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_1
timestamp 1651764895
transform 1 0 1592 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_0_2
timestamp 1651764895
transform 1 0 1608 0 1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_237
timestamp 1651764895
transform 1 0 1624 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_106
timestamp 1651764895
transform 1 0 1672 0 1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_116
timestamp 1651764895
transform -1 0 1784 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_276
timestamp 1651764895
transform 1 0 1784 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_230
timestamp 1651764895
transform 1 0 1848 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_138
timestamp 1651764895
transform 1 0 1912 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_234
timestamp 1651764895
transform -1 0 2040 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_207
timestamp 1651764895
transform 1 0 2040 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_227
timestamp 1651764895
transform 1 0 2072 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_229
timestamp 1651764895
transform 1 0 2136 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_238
timestamp 1651764895
transform 1 0 2184 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_271
timestamp 1651764895
transform 1 0 2232 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_143
timestamp 1651764895
transform 1 0 2296 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_246
timestamp 1651764895
transform -1 0 2392 0 1 3010
box -4 -6 36 206
use NAND2X1  NAND2X1_222
timestamp 1651764895
transform 1 0 2392 0 1 3010
box -4 -6 52 206
use OR2X2  OR2X2_26
timestamp 1651764895
transform 1 0 2440 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_223
timestamp 1651764895
transform -1 0 2552 0 1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_149
timestamp 1651764895
transform -1 0 2616 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_302
timestamp 1651764895
transform -1 0 2680 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_306
timestamp 1651764895
transform 1 0 2680 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_240
timestamp 1651764895
transform 1 0 2744 0 1 3010
box -4 -6 36 206
use AOI21X1  AOI21X1_148
timestamp 1651764895
transform -1 0 2840 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_303
timestamp 1651764895
transform 1 0 2840 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_353
timestamp 1651764895
transform -1 0 2968 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_349
timestamp 1651764895
transform 1 0 2968 0 1 3010
box -4 -6 52 206
use NAND3X1  NAND3X1_310
timestamp 1651764895
transform 1 0 3016 0 1 3010
box -4 -6 68 206
use FILL  FILL_15_1_0
timestamp 1651764895
transform -1 0 3096 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_1
timestamp 1651764895
transform -1 0 3112 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_1_2
timestamp 1651764895
transform -1 0 3128 0 1 3010
box -4 -6 20 206
use OAI21X1  OAI21X1_296
timestamp 1651764895
transform -1 0 3192 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_297
timestamp 1651764895
transform 1 0 3192 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_239
timestamp 1651764895
transform -1 0 3288 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_308
timestamp 1651764895
transform 1 0 3288 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_41
timestamp 1651764895
transform 1 0 3352 0 1 3010
box -4 -6 36 206
use NAND3X1  NAND3X1_399
timestamp 1651764895
transform -1 0 3448 0 1 3010
box -4 -6 68 206
use AND2X2  AND2X2_88
timestamp 1651764895
transform 1 0 3448 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_377
timestamp 1651764895
transform 1 0 3512 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_313
timestamp 1651764895
transform 1 0 3576 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_323
timestamp 1651764895
transform 1 0 3640 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_321
timestamp 1651764895
transform 1 0 3688 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_322
timestamp 1651764895
transform -1 0 3800 0 1 3010
box -4 -6 52 206
use OR2X2  OR2X2_37
timestamp 1651764895
transform -1 0 3864 0 1 3010
box -4 -6 68 206
use NAND2X1  NAND2X1_299
timestamp 1651764895
transform 1 0 3864 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_321
timestamp 1651764895
transform -1 0 3960 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_298
timestamp 1651764895
transform 1 0 3960 0 1 3010
box -4 -6 52 206
use AOI21X1  AOI21X1_152
timestamp 1651764895
transform 1 0 4008 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_314
timestamp 1651764895
transform 1 0 4072 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_315
timestamp 1651764895
transform -1 0 4200 0 1 3010
box -4 -6 68 206
use AOI21X1  AOI21X1_154
timestamp 1651764895
transform 1 0 4200 0 1 3010
box -4 -6 68 206
use INVX1  INVX1_252
timestamp 1651764895
transform 1 0 4264 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_299
timestamp 1651764895
transform -1 0 4360 0 1 3010
box -4 -6 68 206
use NOR3X1  NOR3X1_25
timestamp 1651764895
transform 1 0 4360 0 1 3010
box -4 -6 132 206
use NAND2X1  NAND2X1_363
timestamp 1651764895
transform 1 0 4488 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_373
timestamp 1651764895
transform -1 0 4600 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_169
timestamp 1651764895
transform 1 0 4600 0 1 3010
box -4 -6 52 206
use FILL  FILL_15_2_0
timestamp 1651764895
transform -1 0 4664 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_1
timestamp 1651764895
transform -1 0 4680 0 1 3010
box -4 -6 20 206
use FILL  FILL_15_2_2
timestamp 1651764895
transform -1 0 4696 0 1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_364
timestamp 1651764895
transform -1 0 4744 0 1 3010
box -4 -6 52 206
use NAND2X1  NAND2X1_440
timestamp 1651764895
transform -1 0 4792 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_156
timestamp 1651764895
transform -1 0 4840 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_168
timestamp 1651764895
transform -1 0 4888 0 1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_81
timestamp 1651764895
transform 1 0 4888 0 1 3010
box -4 -6 116 206
use NOR2X1  NOR2X1_133
timestamp 1651764895
transform 1 0 5000 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_134
timestamp 1651764895
transform 1 0 5048 0 1 3010
box -4 -6 52 206
use INVX1  INVX1_266
timestamp 1651764895
transform -1 0 5128 0 1 3010
box -4 -6 36 206
use OAI21X1  OAI21X1_317
timestamp 1651764895
transform -1 0 5192 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_111
timestamp 1651764895
transform 1 0 5192 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_113
timestamp 1651764895
transform 1 0 5240 0 1 3010
box -4 -6 52 206
use NOR2X1  NOR2X1_112
timestamp 1651764895
transform 1 0 5288 0 1 3010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_80
timestamp 1651764895
transform -1 0 5448 0 1 3010
box -4 -6 116 206
use OAI22X1  OAI22X1_8
timestamp 1651764895
transform 1 0 5448 0 1 3010
box -4 -6 84 206
use NAND2X1  NAND2X1_362
timestamp 1651764895
transform -1 0 5576 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_370
timestamp 1651764895
transform -1 0 5640 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_397
timestamp 1651764895
transform -1 0 5704 0 1 3010
box -4 -6 68 206
use NAND3X1  NAND3X1_338
timestamp 1651764895
transform -1 0 5768 0 1 3010
box -4 -6 68 206
use NOR2X1  NOR2X1_131
timestamp 1651764895
transform -1 0 5816 0 1 3010
box -4 -6 52 206
use OAI21X1  OAI21X1_314
timestamp 1651764895
transform 1 0 5816 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_311
timestamp 1651764895
transform -1 0 5944 0 1 3010
box -4 -6 68 206
use OAI21X1  OAI21X1_256
timestamp 1651764895
transform 1 0 5944 0 1 3010
box -4 -6 68 206
use DFFPOSX1  DFFPOSX1_13
timestamp 1651764895
transform 1 0 6008 0 1 3010
box -4 -6 196 206
use BUFX2  BUFX2_30
timestamp 1651764895
transform 1 0 6200 0 1 3010
box -4 -6 52 206
use FILL  FILL_16_1
timestamp 1651764895
transform 1 0 6248 0 1 3010
box -4 -6 20 206
use NAND2X1  NAND2X1_510
timestamp 1651764895
transform 1 0 8 0 -1 3410
box -4 -6 52 206
use XOR2X1  XOR2X1_47
timestamp 1651764895
transform -1 0 168 0 -1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_407
timestamp 1651764895
transform -1 0 216 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_465
timestamp 1651764895
transform -1 0 264 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_344
timestamp 1651764895
transform 1 0 264 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_294
timestamp 1651764895
transform 1 0 312 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_343
timestamp 1651764895
transform -1 0 408 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_245
timestamp 1651764895
transform 1 0 408 0 -1 3410
box -4 -6 36 206
use INVX1  INVX1_179
timestamp 1651764895
transform 1 0 440 0 -1 3410
box -4 -6 36 206
use AND2X2  AND2X2_52
timestamp 1651764895
transform 1 0 472 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_283
timestamp 1651764895
transform 1 0 536 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_282
timestamp 1651764895
transform 1 0 600 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_136
timestamp 1651764895
transform 1 0 664 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_126
timestamp 1651764895
transform -1 0 776 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_293
timestamp 1651764895
transform 1 0 776 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_231
timestamp 1651764895
transform 1 0 824 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_230
timestamp 1651764895
transform 1 0 872 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_229
timestamp 1651764895
transform 1 0 920 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_228
timestamp 1651764895
transform -1 0 1048 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_177
timestamp 1651764895
transform 1 0 1048 0 -1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_122
timestamp 1651764895
transform -1 0 1128 0 -1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_133
timestamp 1651764895
transform -1 0 1192 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_104
timestamp 1651764895
transform -1 0 1240 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_173
timestamp 1651764895
transform 1 0 1240 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_172
timestamp 1651764895
transform 1 0 1288 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_224
timestamp 1651764895
transform 1 0 1336 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_224
timestamp 1651764895
transform 1 0 1384 0 -1 3410
box -4 -6 68 206
use XOR2X1  XOR2X1_13
timestamp 1651764895
transform -1 0 1560 0 -1 3410
box -4 -6 116 206
use FILL  FILL_16_0_0
timestamp 1651764895
transform 1 0 1560 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_1
timestamp 1651764895
transform 1 0 1576 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_0_2
timestamp 1651764895
transform 1 0 1592 0 -1 3410
box -4 -6 20 206
use NOR2X1  NOR2X1_103
timestamp 1651764895
transform 1 0 1608 0 -1 3410
box -4 -6 52 206
use AND2X2  AND2X2_50
timestamp 1651764895
transform 1 0 1656 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_226
timestamp 1651764895
transform 1 0 1720 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_225
timestamp 1651764895
transform 1 0 1784 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_206
timestamp 1651764895
transform -1 0 1880 0 -1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_227
timestamp 1651764895
transform 1 0 1880 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_228
timestamp 1651764895
transform 1 0 1928 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_1
timestamp 1651764895
transform 1 0 1976 0 -1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_226
timestamp 1651764895
transform 1 0 2024 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_233
timestamp 1651764895
transform -1 0 2152 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_284
timestamp 1651764895
transform 1 0 2152 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_289
timestamp 1651764895
transform -1 0 2264 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_291
timestamp 1651764895
transform 1 0 2264 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_298
timestamp 1651764895
transform -1 0 2392 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_296
timestamp 1651764895
transform -1 0 2456 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_297
timestamp 1651764895
transform -1 0 2520 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_147
timestamp 1651764895
transform 1 0 2520 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_301
timestamp 1651764895
transform -1 0 2648 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_300
timestamp 1651764895
transform -1 0 2712 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_293
timestamp 1651764895
transform -1 0 2776 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_292
timestamp 1651764895
transform -1 0 2840 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_274
timestamp 1651764895
transform 1 0 2840 0 -1 3410
box -4 -6 36 206
use AOI21X1  AOI21X1_163
timestamp 1651764895
transform -1 0 2936 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_311
timestamp 1651764895
transform -1 0 3000 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_530
timestamp 1651764895
transform 1 0 3000 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_157
timestamp 1651764895
transform 1 0 3048 0 -1 3410
box -4 -6 52 206
use FILL  FILL_16_1_0
timestamp 1651764895
transform -1 0 3112 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_1
timestamp 1651764895
transform -1 0 3128 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_1_2
timestamp 1651764895
transform -1 0 3144 0 -1 3410
box -4 -6 20 206
use NOR2X1  NOR2X1_172
timestamp 1651764895
transform -1 0 3192 0 -1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_218
timestamp 1651764895
transform -1 0 3256 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_447
timestamp 1651764895
transform -1 0 3304 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_342
timestamp 1651764895
transform -1 0 3336 0 -1 3410
box -4 -6 36 206
use AOI21X1  AOI21X1_219
timestamp 1651764895
transform -1 0 3400 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_309
timestamp 1651764895
transform -1 0 3464 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_426
timestamp 1651764895
transform 1 0 3464 0 -1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_457
timestamp 1651764895
transform -1 0 3592 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_446
timestamp 1651764895
transform 1 0 3592 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_320
timestamp 1651764895
transform 1 0 3640 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_374
timestamp 1651764895
transform 1 0 3688 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_137
timestamp 1651764895
transform 1 0 3736 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_376
timestamp 1651764895
transform -1 0 3848 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_162
timestamp 1651764895
transform -1 0 3912 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_249
timestamp 1651764895
transform -1 0 3944 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_312
timestamp 1651764895
transform -1 0 4008 0 -1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_153
timestamp 1651764895
transform 1 0 4008 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_276
timestamp 1651764895
transform -1 0 4120 0 -1 3410
box -4 -6 52 206
use XOR2X1  XOR2X1_21
timestamp 1651764895
transform -1 0 4232 0 -1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_535
timestamp 1651764895
transform -1 0 4280 0 -1 3410
box -4 -6 52 206
use XOR2X1  XOR2X1_51
timestamp 1651764895
transform -1 0 4392 0 -1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_438
timestamp 1651764895
transform 1 0 4392 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_439
timestamp 1651764895
transform -1 0 4488 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_166
timestamp 1651764895
transform -1 0 4536 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_374
timestamp 1651764895
transform 1 0 4536 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_167
timestamp 1651764895
transform -1 0 4648 0 -1 3410
box -4 -6 52 206
use FILL  FILL_16_2_0
timestamp 1651764895
transform -1 0 4664 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_1
timestamp 1651764895
transform -1 0 4680 0 -1 3410
box -4 -6 20 206
use FILL  FILL_16_2_2
timestamp 1651764895
transform -1 0 4696 0 -1 3410
box -4 -6 20 206
use INVX1  INVX1_334
timestamp 1651764895
transform -1 0 4728 0 -1 3410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_40
timestamp 1651764895
transform 1 0 4728 0 -1 3410
box -4 -6 116 206
use NOR2X1  NOR2X1_132
timestamp 1651764895
transform -1 0 4888 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_110
timestamp 1651764895
transform -1 0 4936 0 -1 3410
box -4 -6 52 206
use INVX1  INVX1_230
timestamp 1651764895
transform 1 0 4936 0 -1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_258
timestamp 1651764895
transform 1 0 4968 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_312
timestamp 1651764895
transform 1 0 5016 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_115
timestamp 1651764895
transform 1 0 5064 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_114
timestamp 1651764895
transform -1 0 5160 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_259
timestamp 1651764895
transform 1 0 5160 0 -1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_199
timestamp 1651764895
transform -1 0 5272 0 -1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_423
timestamp 1651764895
transform 1 0 5272 0 -1 3410
box -4 -6 68 206
use OR2X2  OR2X2_44
timestamp 1651764895
transform 1 0 5336 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_476
timestamp 1651764895
transform -1 0 5464 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_422
timestamp 1651764895
transform -1 0 5528 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_437
timestamp 1651764895
transform 1 0 5528 0 -1 3410
box -4 -6 52 206
use AND2X2  AND2X2_85
timestamp 1651764895
transform 1 0 5576 0 -1 3410
box -4 -6 68 206
use AND2X2  AND2X2_68
timestamp 1651764895
transform 1 0 5640 0 -1 3410
box -4 -6 68 206
use AND2X2  AND2X2_60
timestamp 1651764895
transform -1 0 5768 0 -1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_257
timestamp 1651764895
transform 1 0 5768 0 -1 3410
box -4 -6 68 206
use INVX1  INVX1_228
timestamp 1651764895
transform 1 0 5832 0 -1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_279
timestamp 1651764895
transform -1 0 5928 0 -1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_359
timestamp 1651764895
transform -1 0 5976 0 -1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_491
timestamp 1651764895
transform -1 0 6024 0 -1 3410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_54
timestamp 1651764895
transform 1 0 6024 0 -1 3410
box -4 -6 116 206
use NOR2X1  NOR2X1_153
timestamp 1651764895
transform 1 0 6136 0 -1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_152
timestamp 1651764895
transform -1 0 6232 0 -1 3410
box -4 -6 52 206
use FILL  FILL_17_1
timestamp 1651764895
transform -1 0 6248 0 -1 3410
box -4 -6 20 206
use FILL  FILL_17_2
timestamp 1651764895
transform -1 0 6264 0 -1 3410
box -4 -6 20 206
use XNOR2X1  XNOR2X1_72
timestamp 1651764895
transform 1 0 8 0 1 3410
box -4 -6 116 206
use INVX1  INVX1_319
timestamp 1651764895
transform 1 0 120 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_451
timestamp 1651764895
transform 1 0 152 0 1 3410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_51
timestamp 1651764895
transform 1 0 8 0 -1 3810
box -4 -6 116 206
use OR2X2  OR2X2_56
timestamp 1651764895
transform 1 0 120 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_501
timestamp 1651764895
transform 1 0 184 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_450
timestamp 1651764895
transform -1 0 280 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_397
timestamp 1651764895
transform 1 0 280 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_149
timestamp 1651764895
transform -1 0 392 0 1 3410
box -4 -6 52 206
use INVX1  INVX1_210
timestamp 1651764895
transform 1 0 392 0 1 3410
box -4 -6 36 206
use AND2X2  AND2X2_90
timestamp 1651764895
transform -1 0 296 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_447
timestamp 1651764895
transform 1 0 296 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_188
timestamp 1651764895
transform -1 0 408 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_448
timestamp 1651764895
transform -1 0 472 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_281
timestamp 1651764895
transform -1 0 488 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_159
timestamp 1651764895
transform -1 0 536 0 1 3410
box -4 -6 52 206
use OAI22X1  OAI22X1_9
timestamp 1651764895
transform 1 0 536 0 1 3410
box -4 -6 84 206
use NAND2X1  NAND2X1_406
timestamp 1651764895
transform -1 0 520 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_342
timestamp 1651764895
transform -1 0 568 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_340
timestamp 1651764895
transform 1 0 568 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_244
timestamp 1651764895
transform 1 0 616 0 1 3410
box -4 -6 36 206
use AOI21X1  AOI21X1_170
timestamp 1651764895
transform 1 0 648 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_280
timestamp 1651764895
transform 1 0 712 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_340
timestamp 1651764895
transform 1 0 776 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_290
timestamp 1651764895
transform 1 0 616 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_339
timestamp 1651764895
transform -1 0 728 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_148
timestamp 1651764895
transform 1 0 728 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_75
timestamp 1651764895
transform 1 0 776 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_135
timestamp 1651764895
transform 1 0 840 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_287
timestamp 1651764895
transform 1 0 904 0 1 3410
box -4 -6 68 206
use NOR3X1  NOR3X1_23
timestamp 1651764895
transform -1 0 1096 0 1 3410
box -4 -6 132 206
use OAI21X1  OAI21X1_277
timestamp 1651764895
transform 1 0 840 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_232
timestamp 1651764895
transform 1 0 904 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_278
timestamp 1651764895
transform 1 0 952 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_286
timestamp 1651764895
transform 1 0 1096 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_284
timestamp 1651764895
transform 1 0 1160 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_146
timestamp 1651764895
transform -1 0 1064 0 -1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_168
timestamp 1651764895
transform -1 0 1128 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_45
timestamp 1651764895
transform 1 0 1128 0 -1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_124
timestamp 1651764895
transform -1 0 1208 0 -1 3810
box -4 -6 52 206
use XOR2X1  XOR2X1_20
timestamp 1651764895
transform 1 0 1208 0 -1 3810
box -4 -6 116 206
use NAND3X1  NAND3X1_291
timestamp 1651764895
transform 1 0 1224 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_137
timestamp 1651764895
transform 1 0 1288 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_288
timestamp 1651764895
transform 1 0 1352 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_337
timestamp 1651764895
transform 1 0 1320 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_225
timestamp 1651764895
transform 1 0 1384 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_272
timestamp 1651764895
transform 1 0 1480 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_226
timestamp 1651764895
transform 1 0 1432 0 -1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_139
timestamp 1651764895
transform 1 0 1480 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_223
timestamp 1651764895
transform 1 0 1416 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_285
timestamp 1651764895
transform 1 0 1544 0 -1 3810
box -4 -6 52 206
use FILL  FILL_17_0_0
timestamp 1651764895
transform 1 0 1544 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_0_1
timestamp 1651764895
transform -1 0 1624 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_0_0
timestamp 1651764895
transform -1 0 1608 0 -1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_285
timestamp 1651764895
transform 1 0 1592 0 1 3410
box -4 -6 68 206
use FILL  FILL_17_0_2
timestamp 1651764895
transform 1 0 1576 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_0_1
timestamp 1651764895
transform 1 0 1560 0 1 3410
box -4 -6 20 206
use AOI21X1  AOI21X1_173
timestamp 1651764895
transform -1 0 1720 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_140
timestamp 1651764895
transform 1 0 1720 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_289
timestamp 1651764895
transform 1 0 1784 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_0_2
timestamp 1651764895
transform -1 0 1640 0 -1 3810
box -4 -6 20 206
use XNOR2X1  XNOR2X1_34
timestamp 1651764895
transform -1 0 1752 0 -1 3810
box -4 -6 116 206
use OAI21X1  OAI21X1_273
timestamp 1651764895
transform -1 0 1816 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_120
timestamp 1651764895
transform 1 0 1848 0 1 3410
box -4 -6 52 206
use NOR3X1  NOR3X1_24
timestamp 1651764895
transform -1 0 2024 0 1 3410
box -4 -6 132 206
use NOR2X1  NOR2X1_123
timestamp 1651764895
transform -1 0 1864 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_62
timestamp 1651764895
transform 1 0 1864 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_274
timestamp 1651764895
transform 1 0 1928 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_275
timestamp 1651764895
transform 1 0 1992 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_287
timestamp 1651764895
transform 1 0 2024 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_288
timestamp 1651764895
transform 1 0 2088 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_294
timestamp 1651764895
transform -1 0 2216 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_243
timestamp 1651764895
transform 1 0 2056 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_288
timestamp 1651764895
transform 1 0 2088 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_287
timestamp 1651764895
transform 1 0 2136 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_73
timestamp 1651764895
transform 1 0 2184 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_142
timestamp 1651764895
transform 1 0 2216 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_144
timestamp 1651764895
transform 1 0 2280 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_290
timestamp 1651764895
transform 1 0 2344 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_121
timestamp 1651764895
transform 1 0 2408 0 1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_286
timestamp 1651764895
transform -1 0 2312 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_293
timestamp 1651764895
transform -1 0 2376 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_176
timestamp 1651764895
transform -1 0 2440 0 -1 3810
box -4 -6 68 206
use OR2X2  OR2X2_29
timestamp 1651764895
transform 1 0 2456 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_290
timestamp 1651764895
transform 1 0 2520 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_295
timestamp 1651764895
transform -1 0 2632 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_289
timestamp 1651764895
transform -1 0 2488 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_285
timestamp 1651764895
transform 1 0 2488 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_292
timestamp 1651764895
transform 1 0 2552 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_331
timestamp 1651764895
transform 1 0 2632 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_141
timestamp 1651764895
transform -1 0 2760 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_295
timestamp 1651764895
transform 1 0 2760 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_331
timestamp 1651764895
transform -1 0 2664 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_289
timestamp 1651764895
transform 1 0 2664 0 -1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_179
timestamp 1651764895
transform -1 0 2760 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_330
timestamp 1651764895
transform 1 0 2760 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_275
timestamp 1651764895
transform -1 0 2840 0 -1 3810
box -4 -6 36 206
use XOR2X1  XOR2X1_18
timestamp 1651764895
transform -1 0 2936 0 1 3410
box -4 -6 116 206
use AOI21X1  AOI21X1_146
timestamp 1651764895
transform -1 0 3000 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_299
timestamp 1651764895
transform 1 0 3000 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_348
timestamp 1651764895
transform 1 0 2840 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_352
timestamp 1651764895
transform 1 0 2888 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1651764895
transform 1 0 2936 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_353
timestamp 1651764895
transform 1 0 2968 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_501
timestamp 1651764895
transform 1 0 3064 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_7
timestamp 1651764895
transform 1 0 3016 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_367
timestamp 1651764895
transform 1 0 3064 0 1 3410
box -4 -6 68 206
use FILL  FILL_18_1_2
timestamp 1651764895
transform -1 0 3176 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_1
timestamp 1651764895
transform -1 0 3160 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_1_0
timestamp 1651764895
transform -1 0 3144 0 -1 3810
box -4 -6 20 206
use FILL  FILL_17_1_2
timestamp 1651764895
transform -1 0 3176 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_1
timestamp 1651764895
transform -1 0 3160 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_1_0
timestamp 1651764895
transform -1 0 3144 0 1 3410
box -4 -6 20 206
use NOR2X1  NOR2X1_196
timestamp 1651764895
transform -1 0 3224 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_6
timestamp 1651764895
transform -1 0 3224 0 1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_525
timestamp 1651764895
transform -1 0 3288 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_500
timestamp 1651764895
transform -1 0 3352 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_8
timestamp 1651764895
transform -1 0 3400 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_9
timestamp 1651764895
transform 1 0 3400 0 1 3410
box -4 -6 52 206
use AOI21X1  AOI21X1_254
timestamp 1651764895
transform -1 0 3288 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_531
timestamp 1651764895
transform -1 0 3336 0 -1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_198
timestamp 1651764895
transform -1 0 3384 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_532
timestamp 1651764895
transform -1 0 3432 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_499
timestamp 1651764895
transform 1 0 3448 0 1 3410
box -4 -6 68 206
use NOR2X1  NOR2X1_197
timestamp 1651764895
transform 1 0 3512 0 1 3410
box -4 -6 52 206
use NAND2X1  NAND2X1_297
timestamp 1651764895
transform 1 0 3560 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_498
timestamp 1651764895
transform -1 0 3672 0 1 3410
box -4 -6 68 206
use AOI21X1  AOI21X1_185
timestamp 1651764895
transform -1 0 3496 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_329
timestamp 1651764895
transform -1 0 3544 0 -1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_196
timestamp 1651764895
transform 1 0 3544 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1651764895
transform 1 0 3608 0 -1 3810
box -4 -6 36 206
use INVX1  INVX1_343
timestamp 1651764895
transform 1 0 3672 0 1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_458
timestamp 1651764895
transform -1 0 3768 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_344
timestamp 1651764895
transform 1 0 3768 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_427
timestamp 1651764895
transform -1 0 3864 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_273
timestamp 1651764895
transform -1 0 3672 0 -1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_138
timestamp 1651764895
transform -1 0 3720 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_448
timestamp 1651764895
transform -1 0 3768 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_100
timestamp 1651764895
transform 1 0 3768 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_345
timestamp 1651764895
transform 1 0 3864 0 1 3410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_38
timestamp 1651764895
transform 1 0 3896 0 1 3410
box -4 -6 116 206
use XOR2X1  XOR2X1_22
timestamp 1651764895
transform -1 0 4120 0 1 3410
box -4 -6 116 206
use XNOR2X1  XNOR2X1_43
timestamp 1651764895
transform 1 0 3832 0 -1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_324
timestamp 1651764895
transform 1 0 3944 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_375
timestamp 1651764895
transform 1 0 3992 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_325
timestamp 1651764895
transform 1 0 4120 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_322
timestamp 1651764895
transform -1 0 4232 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_375
timestamp 1651764895
transform 1 0 4056 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_342
timestamp 1651764895
transform -1 0 4184 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_328
timestamp 1651764895
transform -1 0 4232 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_327
timestamp 1651764895
transform 1 0 4232 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_323
timestamp 1651764895
transform 1 0 4280 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_272
timestamp 1651764895
transform 1 0 4344 0 1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_343
timestamp 1651764895
transform 1 0 4376 0 1 3410
box -4 -6 68 206
use AND2X2  AND2X2_80
timestamp 1651764895
transform 1 0 4232 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_326
timestamp 1651764895
transform 1 0 4296 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_87
timestamp 1651764895
transform 1 0 4344 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_355
timestamp 1651764895
transform 1 0 4408 0 -1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_376
timestamp 1651764895
transform 1 0 4440 0 1 3410
box -4 -6 68 206
use OR2X2  OR2X2_45
timestamp 1651764895
transform -1 0 4568 0 1 3410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_78
timestamp 1651764895
transform 1 0 4568 0 1 3410
box -4 -6 116 206
use INVX1  INVX1_335
timestamp 1651764895
transform -1 0 4488 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_441
timestamp 1651764895
transform -1 0 4536 0 -1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_424
timestamp 1651764895
transform -1 0 4600 0 -1 3810
box -4 -6 68 206
use AND2X2  AND2X2_71
timestamp 1651764895
transform -1 0 4664 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_2_1
timestamp 1651764895
transform -1 0 4696 0 -1 3810
box -4 -6 20 206
use FILL  FILL_18_2_0
timestamp 1651764895
transform -1 0 4680 0 -1 3810
box -4 -6 20 206
use FILL  FILL_17_2_0
timestamp 1651764895
transform 1 0 4680 0 1 3410
box -4 -6 20 206
use OAI21X1  OAI21X1_318
timestamp 1651764895
transform 1 0 4760 0 -1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_135
timestamp 1651764895
transform -1 0 4760 0 -1 3810
box -4 -6 52 206
use FILL  FILL_18_2_2
timestamp 1651764895
transform -1 0 4712 0 -1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_506
timestamp 1651764895
transform -1 0 4824 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_338
timestamp 1651764895
transform 1 0 4728 0 1 3410
box -4 -6 36 206
use FILL  FILL_17_2_2
timestamp 1651764895
transform 1 0 4712 0 1 3410
box -4 -6 20 206
use FILL  FILL_17_2_1
timestamp 1651764895
transform 1 0 4696 0 1 3410
box -4 -6 20 206
use NAND2X1  NAND2X1_314
timestamp 1651764895
transform 1 0 4856 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_267
timestamp 1651764895
transform -1 0 4856 0 -1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_455
timestamp 1651764895
transform 1 0 4888 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_336
timestamp 1651764895
transform -1 0 4888 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_337
timestamp 1651764895
transform -1 0 4856 0 1 3410
box -4 -6 36 206
use NAND2X1  NAND2X1_316
timestamp 1651764895
transform 1 0 4952 0 -1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_318
timestamp 1651764895
transform -1 0 4952 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_70
timestamp 1651764895
transform -1 0 5016 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_317
timestamp 1651764895
transform -1 0 5048 0 -1 3810
box -4 -6 52 206
use OR2X2  OR2X2_30
timestamp 1651764895
transform -1 0 5080 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_372
timestamp 1651764895
transform -1 0 5144 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_316
timestamp 1651764895
transform 1 0 5144 0 1 3410
box -4 -6 68 206
use NAND3X1  NAND3X1_280
timestamp 1651764895
transform -1 0 5272 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_268
timestamp 1651764895
transform 1 0 5048 0 -1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_315
timestamp 1651764895
transform -1 0 5128 0 -1 3810
box -4 -6 52 206
use AND2X2  AND2X2_86
timestamp 1651764895
transform -1 0 5192 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_371
timestamp 1651764895
transform -1 0 5256 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_129
timestamp 1651764895
transform 1 0 5272 0 1 3410
box -4 -6 68 206
use AND2X2  AND2X2_98
timestamp 1651764895
transform -1 0 5400 0 1 3410
box -4 -6 68 206
use OAI21X1  OAI21X1_313
timestamp 1651764895
transform -1 0 5464 0 1 3410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_56
timestamp 1651764895
transform 1 0 5256 0 -1 3810
box -4 -6 116 206
use AND2X2  AND2X2_97
timestamp 1651764895
transform -1 0 5432 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_231
timestamp 1651764895
transform 1 0 5464 0 1 3410
box -4 -6 36 206
use NOR2X1  NOR2X1_116
timestamp 1651764895
transform -1 0 5544 0 1 3410
box -4 -6 52 206
use OAI21X1  OAI21X1_260
timestamp 1651764895
transform 1 0 5544 0 1 3410
box -4 -6 68 206
use NAND2X1  NAND2X1_260
timestamp 1651764895
transform 1 0 5608 0 1 3410
box -4 -6 52 206
use AND2X2  AND2X2_82
timestamp 1651764895
transform -1 0 5496 0 -1 3810
box -4 -6 68 206
use AND2X2  AND2X2_69
timestamp 1651764895
transform -1 0 5560 0 -1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_315
timestamp 1651764895
transform 1 0 5560 0 -1 3810
box -4 -6 68 206
use INVX1  INVX1_299
timestamp 1651764895
transform -1 0 5720 0 -1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_419
timestamp 1651764895
transform 1 0 5624 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_259
timestamp 1651764895
transform -1 0 5704 0 1 3410
box -4 -6 52 206
use NOR2X1  NOR2X1_154
timestamp 1651764895
transform -1 0 5800 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_259
timestamp 1651764895
transform -1 0 5752 0 -1 3810
box -4 -6 36 206
use INVX1  INVX1_304
timestamp 1651764895
transform -1 0 5768 0 1 3410
box -4 -6 36 206
use INVX1  INVX1_232
timestamp 1651764895
transform -1 0 5736 0 1 3410
box -4 -6 36 206
use OAI21X1  OAI21X1_367
timestamp 1651764895
transform 1 0 5800 0 -1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_398
timestamp 1651764895
transform -1 0 5864 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_265
timestamp 1651764895
transform -1 0 5800 0 1 3410
box -4 -6 36 206
use NAND3X1  NAND3X1_339
timestamp 1651764895
transform -1 0 5928 0 1 3410
box -4 -6 68 206
use INVX1  INVX1_226
timestamp 1651764895
transform -1 0 5960 0 1 3410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_55
timestamp 1651764895
transform 1 0 5960 0 1 3410
box -4 -6 116 206
use INVX1  INVX1_298
timestamp 1651764895
transform -1 0 5896 0 -1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_393
timestamp 1651764895
transform -1 0 5960 0 -1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_428
timestamp 1651764895
transform -1 0 6008 0 -1 3810
box -4 -6 52 206
use INVX1  INVX1_297
timestamp 1651764895
transform 1 0 6008 0 -1 3810
box -4 -6 36 206
use XOR2X1  XOR2X1_41
timestamp 1651764895
transform 1 0 6072 0 1 3410
box -4 -6 116 206
use NAND2X1  NAND2X1_356
timestamp 1651764895
transform 1 0 6184 0 1 3410
box -4 -6 52 206
use NAND3X1  NAND3X1_396
timestamp 1651764895
transform 1 0 6040 0 -1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_194
timestamp 1651764895
transform -1 0 6168 0 -1 3810
box -4 -6 68 206
use OR2X2  OR2X2_42
timestamp 1651764895
transform -1 0 6232 0 -1 3810
box -4 -6 68 206
use FILL  FILL_18_1
timestamp 1651764895
transform 1 0 6232 0 1 3410
box -4 -6 20 206
use FILL  FILL_18_2
timestamp 1651764895
transform 1 0 6248 0 1 3410
box -4 -6 20 206
use FILL  FILL_19_1
timestamp 1651764895
transform -1 0 6248 0 -1 3810
box -4 -6 20 206
use FILL  FILL_19_2
timestamp 1651764895
transform -1 0 6264 0 -1 3810
box -4 -6 20 206
use XOR2X1  XOR2X1_37
timestamp 1651764895
transform 1 0 8 0 1 3810
box -4 -6 116 206
use OAI21X1  OAI21X1_489
timestamp 1651764895
transform -1 0 184 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_511
timestamp 1651764895
transform -1 0 248 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_160
timestamp 1651764895
transform -1 0 296 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_40
timestamp 1651764895
transform 1 0 296 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_449
timestamp 1651764895
transform -1 0 424 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_396
timestamp 1651764895
transform 1 0 424 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_318
timestamp 1651764895
transform -1 0 520 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_410
timestamp 1651764895
transform 1 0 520 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_462
timestamp 1651764895
transform 1 0 584 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_285
timestamp 1651764895
transform 1 0 632 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_353
timestamp 1651764895
transform 1 0 664 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_286
timestamp 1651764895
transform -1 0 760 0 1 3810
box -4 -6 36 206
use OAI21X1  OAI21X1_393
timestamp 1651764895
transform -1 0 824 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_338
timestamp 1651764895
transform 1 0 824 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_444
timestamp 1651764895
transform 1 0 888 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_443
timestamp 1651764895
transform 1 0 952 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_397
timestamp 1651764895
transform 1 0 1016 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_445
timestamp 1651764895
transform -1 0 1128 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_337
timestamp 1651764895
transform 1 0 1128 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_392
timestamp 1651764895
transform 1 0 1176 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_391
timestamp 1651764895
transform -1 0 1304 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_332
timestamp 1651764895
transform 1 0 1304 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_286
timestamp 1651764895
transform 1 0 1368 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_146
timestamp 1651764895
transform 1 0 1416 0 1 3810
box -4 -6 36 206
use OR2X2  OR2X2_32
timestamp 1651764895
transform 1 0 1448 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_167
timestamp 1651764895
transform 1 0 1512 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_0_0
timestamp 1651764895
transform 1 0 1576 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_1
timestamp 1651764895
transform 1 0 1592 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_0_2
timestamp 1651764895
transform 1 0 1608 0 1 3810
box -4 -6 20 206
use NOR2X1  NOR2X1_144
timestamp 1651764895
transform 1 0 1624 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_283
timestamp 1651764895
transform 1 0 1672 0 1 3810
box -4 -6 36 206
use XOR2X1  XOR2X1_19
timestamp 1651764895
transform -1 0 1816 0 1 3810
box -4 -6 116 206
use NOR2X1  NOR2X1_142
timestamp 1651764895
transform -1 0 1864 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_34
timestamp 1651764895
transform 1 0 1864 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_143
timestamp 1651764895
transform 1 0 1928 0 1 3810
box -4 -6 52 206
use NOR3X1  NOR3X1_26
timestamp 1651764895
transform -1 0 2104 0 1 3810
box -4 -6 132 206
use OAI21X1  OAI21X1_336
timestamp 1651764895
transform 1 0 2104 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_352
timestamp 1651764895
transform 1 0 2168 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_166
timestamp 1651764895
transform -1 0 2296 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_328
timestamp 1651764895
transform -1 0 2360 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_281
timestamp 1651764895
transform -1 0 2392 0 1 3810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_35
timestamp 1651764895
transform 1 0 2392 0 1 3810
box -4 -6 116 206
use AND2X2  AND2X2_79
timestamp 1651764895
transform -1 0 2568 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_346
timestamp 1651764895
transform 1 0 2568 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_406
timestamp 1651764895
transform -1 0 2680 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_291
timestamp 1651764895
transform -1 0 2712 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_350
timestamp 1651764895
transform 1 0 2712 0 1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_477
timestamp 1651764895
transform 1 0 2760 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_351
timestamp 1651764895
transform 1 0 2824 0 1 3810
box -4 -6 52 206
use AOI21X1  AOI21X1_211
timestamp 1651764895
transform 1 0 2872 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_526
timestamp 1651764895
transform -1 0 3000 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_378
timestamp 1651764895
transform 1 0 3000 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_530
timestamp 1651764895
transform 1 0 3032 0 1 3810
box -4 -6 68 206
use FILL  FILL_19_1_0
timestamp 1651764895
transform -1 0 3112 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_1
timestamp 1651764895
transform -1 0 3128 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_1_2
timestamp 1651764895
transform -1 0 3144 0 1 3810
box -4 -6 20 206
use OAI21X1  OAI21X1_502
timestamp 1651764895
transform -1 0 3208 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_174
timestamp 1651764895
transform 1 0 3208 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_504
timestamp 1651764895
transform 1 0 3256 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_355
timestamp 1651764895
transform 1 0 3320 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_369
timestamp 1651764895
transform -1 0 3448 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_366
timestamp 1651764895
transform -1 0 3512 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_356
timestamp 1651764895
transform -1 0 3576 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_187
timestamp 1651764895
transform 1 0 3576 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_368
timestamp 1651764895
transform 1 0 3640 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_370
timestamp 1651764895
transform -1 0 3768 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_186
timestamp 1651764895
transform 1 0 3768 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_359
timestamp 1651764895
transform 1 0 3832 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_358
timestamp 1651764895
transform 1 0 3896 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_373
timestamp 1651764895
transform -1 0 4024 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_378
timestamp 1651764895
transform -1 0 4088 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_374
timestamp 1651764895
transform 1 0 4088 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_372
timestamp 1651764895
transform 1 0 4152 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_377
timestamp 1651764895
transform 1 0 4216 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_379
timestamp 1651764895
transform -1 0 4344 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_189
timestamp 1651764895
transform 1 0 4344 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_381
timestamp 1651764895
transform -1 0 4472 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_333
timestamp 1651764895
transform -1 0 4504 0 1 3810
box -4 -6 36 206
use AOI21X1  AOI21X1_195
timestamp 1651764895
transform 1 0 4504 0 1 3810
box -4 -6 68 206
use NOR2X1  NOR2X1_136
timestamp 1651764895
transform -1 0 4616 0 1 3810
box -4 -6 52 206
use NAND2X1  NAND2X1_313
timestamp 1651764895
transform -1 0 4664 0 1 3810
box -4 -6 52 206
use FILL  FILL_19_2_0
timestamp 1651764895
transform 1 0 4664 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_1
timestamp 1651764895
transform 1 0 4680 0 1 3810
box -4 -6 20 206
use FILL  FILL_19_2_2
timestamp 1651764895
transform 1 0 4696 0 1 3810
box -4 -6 20 206
use XNOR2X1  XNOR2X1_41
timestamp 1651764895
transform 1 0 4712 0 1 3810
box -4 -6 116 206
use NAND2X1  NAND2X1_435
timestamp 1651764895
transform -1 0 4872 0 1 3810
box -4 -6 52 206
use NAND3X1  NAND3X1_341
timestamp 1651764895
transform -1 0 4936 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_269
timestamp 1651764895
transform -1 0 4968 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_340
timestamp 1651764895
transform -1 0 5032 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_305
timestamp 1651764895
transform -1 0 5064 0 1 3810
box -4 -6 36 206
use INVX1  INVX1_365
timestamp 1651764895
transform 1 0 5064 0 1 3810
box -4 -6 36 206
use NOR2X1  NOR2X1_165
timestamp 1651764895
transform 1 0 5096 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_474
timestamp 1651764895
transform 1 0 5144 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_430
timestamp 1651764895
transform -1 0 5256 0 1 3810
box -4 -6 52 206
use OR2X2  OR2X2_43
timestamp 1651764895
transform -1 0 5320 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_429
timestamp 1651764895
transform -1 0 5368 0 1 3810
box -4 -6 52 206
use NOR2X1  NOR2X1_164
timestamp 1651764895
transform 1 0 5368 0 1 3810
box -4 -6 52 206
use XOR2X1  XOR2X1_25
timestamp 1651764895
transform 1 0 5416 0 1 3810
box -4 -6 116 206
use NOR2X1  NOR2X1_163
timestamp 1651764895
transform 1 0 5528 0 1 3810
box -4 -6 52 206
use OAI21X1  OAI21X1_312
timestamp 1651764895
transform -1 0 5640 0 1 3810
box -4 -6 68 206
use OAI21X1  OAI21X1_368
timestamp 1651764895
transform 1 0 5640 0 1 3810
box -4 -6 68 206
use NAND2X1  NAND2X1_306
timestamp 1651764895
transform -1 0 5752 0 1 3810
box -4 -6 52 206
use INVX1  INVX1_260
timestamp 1651764895
transform -1 0 5784 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_395
timestamp 1651764895
transform -1 0 5848 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_392
timestamp 1651764895
transform -1 0 5912 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_258
timestamp 1651764895
transform -1 0 5944 0 1 3810
box -4 -6 36 206
use NAND3X1  NAND3X1_390
timestamp 1651764895
transform 1 0 5944 0 1 3810
box -4 -6 68 206
use NAND3X1  NAND3X1_394
timestamp 1651764895
transform -1 0 6072 0 1 3810
box -4 -6 68 206
use AOI21X1  AOI21X1_193
timestamp 1651764895
transform 1 0 6072 0 1 3810
box -4 -6 68 206
use INVX1  INVX1_296
timestamp 1651764895
transform -1 0 6168 0 1 3810
box -4 -6 36 206
use NAND2X1  NAND2X1_425
timestamp 1651764895
transform -1 0 6216 0 1 3810
box -4 -6 52 206
use FILL  FILL_20_1
timestamp 1651764895
transform 1 0 6216 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_2
timestamp 1651764895
transform 1 0 6232 0 1 3810
box -4 -6 20 206
use FILL  FILL_20_3
timestamp 1651764895
transform 1 0 6248 0 1 3810
box -4 -6 20 206
use XNOR2X1  XNOR2X1_69
timestamp 1651764895
transform 1 0 8 0 -1 4210
box -4 -6 116 206
use XOR2X1  XOR2X1_48
timestamp 1651764895
transform 1 0 120 0 -1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_507
timestamp 1651764895
transform -1 0 280 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_485
timestamp 1651764895
transform -1 0 344 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_405
timestamp 1651764895
transform 1 0 344 0 -1 4210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_52
timestamp 1651764895
transform -1 0 504 0 -1 4210
box -4 -6 116 206
use NOR3X1  NOR3X1_27
timestamp 1651764895
transform -1 0 632 0 -1 4210
box -4 -6 132 206
use OAI21X1  OAI21X1_341
timestamp 1651764895
transform 1 0 632 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_463
timestamp 1651764895
transform -1 0 744 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_51
timestamp 1651764895
transform -1 0 808 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_396
timestamp 1651764895
transform -1 0 856 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_343
timestamp 1651764895
transform 1 0 856 0 -1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_28
timestamp 1651764895
transform 1 0 920 0 -1 4210
box -4 -6 132 206
use NAND2X1  NAND2X1_341
timestamp 1651764895
transform -1 0 1096 0 -1 4210
box -4 -6 52 206
use AND2X2  AND2X2_77
timestamp 1651764895
transform 1 0 1096 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_339
timestamp 1651764895
transform 1 0 1160 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_442
timestamp 1651764895
transform 1 0 1208 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_333
timestamp 1651764895
transform 1 0 1272 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_50
timestamp 1651764895
transform -1 0 1368 0 -1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_395
timestamp 1651764895
transform 1 0 1368 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_394
timestamp 1651764895
transform 1 0 1416 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_399
timestamp 1651764895
transform 1 0 1480 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_39
timestamp 1651764895
transform -1 0 1592 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_0_0
timestamp 1651764895
transform -1 0 1608 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_1
timestamp 1651764895
transform -1 0 1624 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_0_2
timestamp 1651764895
transform -1 0 1640 0 -1 4210
box -4 -6 20 206
use OAI21X1  OAI21X1_390
timestamp 1651764895
transform -1 0 1704 0 -1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_28
timestamp 1651764895
transform -1 0 1816 0 -1 4210
box -4 -6 116 206
use OAI21X1  OAI21X1_334
timestamp 1651764895
transform 1 0 1816 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_145
timestamp 1651764895
transform 1 0 1880 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_33
timestamp 1651764895
transform 1 0 1928 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_335
timestamp 1651764895
transform -1 0 2056 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_386
timestamp 1651764895
transform 1 0 2056 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_284
timestamp 1651764895
transform 1 0 2120 0 -1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_169
timestamp 1651764895
transform -1 0 2216 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_351
timestamp 1651764895
transform 1 0 2216 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_349
timestamp 1651764895
transform 1 0 2280 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_182
timestamp 1651764895
transform 1 0 2344 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_348
timestamp 1651764895
transform 1 0 2408 0 -1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_34
timestamp 1651764895
transform -1 0 2600 0 -1 4210
box -4 -6 132 206
use OAI21X1  OAI21X1_352
timestamp 1651764895
transform 1 0 2600 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_365
timestamp 1651764895
transform 1 0 2664 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_351
timestamp 1651764895
transform 1 0 2728 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_479
timestamp 1651764895
transform 1 0 2792 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_412
timestamp 1651764895
transform 1 0 2856 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_410
timestamp 1651764895
transform -1 0 2952 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_427
timestamp 1651764895
transform 1 0 2952 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_5
timestamp 1651764895
transform 1 0 3016 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_527
timestamp 1651764895
transform 1 0 3064 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_1_0
timestamp 1651764895
transform 1 0 3128 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_1
timestamp 1651764895
transform 1 0 3144 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_1_2
timestamp 1651764895
transform 1 0 3160 0 -1 4210
box -4 -6 20 206
use NAND2X1  NAND2X1_411
timestamp 1651764895
transform 1 0 3176 0 -1 4210
box -4 -6 52 206
use AOI21X1  AOI21X1_228
timestamp 1651764895
transform 1 0 3224 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_432
timestamp 1651764895
transform -1 0 3352 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_428
timestamp 1651764895
transform -1 0 3416 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_375
timestamp 1651764895
transform 1 0 3416 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_414
timestamp 1651764895
transform 1 0 3464 0 -1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_173
timestamp 1651764895
transform -1 0 3560 0 -1 4210
box -4 -6 52 206
use AOI22X1  AOI22X1_45
timestamp 1651764895
transform -1 0 3640 0 -1 4210
box -4 -6 84 206
use OAI21X1  OAI21X1_428
timestamp 1651764895
transform 1 0 3640 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_450
timestamp 1651764895
transform 1 0 3704 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_378
timestamp 1651764895
transform 1 0 3752 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_449
timestamp 1651764895
transform 1 0 3816 0 -1 4210
box -4 -6 52 206
use XOR2X1  XOR2X1_26
timestamp 1651764895
transform 1 0 3864 0 -1 4210
box -4 -6 116 206
use AND2X2  AND2X2_89
timestamp 1651764895
transform 1 0 3976 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_294
timestamp 1651764895
transform -1 0 4072 0 -1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_371
timestamp 1651764895
transform -1 0 4136 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_381
timestamp 1651764895
transform -1 0 4184 0 -1 4210
box -4 -6 52 206
use OR2X2  OR2X2_59
timestamp 1651764895
transform -1 0 4248 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_537
timestamp 1651764895
transform -1 0 4296 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_380
timestamp 1651764895
transform -1 0 4360 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_188
timestamp 1651764895
transform -1 0 4424 0 -1 4210
box -4 -6 68 206
use OR2X2  OR2X2_46
timestamp 1651764895
transform -1 0 4488 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_442
timestamp 1651764895
transform -1 0 4536 0 -1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_369
timestamp 1651764895
transform -1 0 4584 0 -1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_383
timestamp 1651764895
transform 1 0 4584 0 -1 4210
box -4 -6 68 206
use FILL  FILL_20_2_0
timestamp 1651764895
transform 1 0 4648 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_1
timestamp 1651764895
transform 1 0 4664 0 -1 4210
box -4 -6 20 206
use FILL  FILL_20_2_2
timestamp 1651764895
transform 1 0 4680 0 -1 4210
box -4 -6 20 206
use INVX1  INVX1_271
timestamp 1651764895
transform 1 0 4696 0 -1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_360
timestamp 1651764895
transform -1 0 4792 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_361
timestamp 1651764895
transform 1 0 4792 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_421
timestamp 1651764895
transform -1 0 4920 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_382
timestamp 1651764895
transform -1 0 4984 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_191
timestamp 1651764895
transform 1 0 4984 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_319
timestamp 1651764895
transform -1 0 5096 0 -1 4210
box -4 -6 52 206
use AOI22X1  AOI22X1_42
timestamp 1651764895
transform 1 0 5096 0 -1 4210
box -4 -6 84 206
use AND2X2  AND2X2_84
timestamp 1651764895
transform 1 0 5176 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_362
timestamp 1651764895
transform 1 0 5240 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_363
timestamp 1651764895
transform 1 0 5304 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_385
timestamp 1651764895
transform -1 0 5432 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_387
timestamp 1651764895
transform 1 0 5432 0 -1 4210
box -4 -6 68 206
use NOR2X1  NOR2X1_130
timestamp 1651764895
transform -1 0 5544 0 -1 4210
box -4 -6 52 206
use INVX1  INVX1_261
timestamp 1651764895
transform 1 0 5544 0 -1 4210
box -4 -6 36 206
use AND2X2  AND2X2_66
timestamp 1651764895
transform 1 0 5576 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_388
timestamp 1651764895
transform -1 0 5704 0 -1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_192
timestamp 1651764895
transform 1 0 5704 0 -1 4210
box -4 -6 68 206
use INVX1  INVX1_264
timestamp 1651764895
transform 1 0 5768 0 -1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_386
timestamp 1651764895
transform 1 0 5800 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_391
timestamp 1651764895
transform 1 0 5864 0 -1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_389
timestamp 1651764895
transform -1 0 5992 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_365
timestamp 1651764895
transform -1 0 6056 0 -1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_364
timestamp 1651764895
transform 1 0 6056 0 -1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_490
timestamp 1651764895
transform -1 0 6168 0 -1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_420
timestamp 1651764895
transform 1 0 6168 0 -1 4210
box -4 -6 68 206
use FILL  FILL_21_1
timestamp 1651764895
transform -1 0 6248 0 -1 4210
box -4 -6 20 206
use FILL  FILL_21_2
timestamp 1651764895
transform -1 0 6264 0 -1 4210
box -4 -6 20 206
use NAND2X1  NAND2X1_466
timestamp 1651764895
transform 1 0 8 0 1 4210
box -4 -6 52 206
use OR2X2  OR2X2_52
timestamp 1651764895
transform -1 0 120 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_487
timestamp 1651764895
transform 1 0 120 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_513
timestamp 1651764895
transform -1 0 248 0 1 4210
box -4 -6 68 206
use OR2X2  OR2X2_57
timestamp 1651764895
transform -1 0 312 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_467
timestamp 1651764895
transform -1 0 360 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_288
timestamp 1651764895
transform 1 0 360 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_354
timestamp 1651764895
transform -1 0 456 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_171
timestamp 1651764895
transform 1 0 456 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_287
timestamp 1651764895
transform -1 0 552 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_408
timestamp 1651764895
transform 1 0 552 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_395
timestamp 1651764895
transform -1 0 664 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_412
timestamp 1651764895
transform -1 0 728 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_172
timestamp 1651764895
transform 1 0 728 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_355
timestamp 1651764895
transform 1 0 792 0 1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_29
timestamp 1651764895
transform -1 0 984 0 1 4210
box -4 -6 132 206
use OAI21X1  OAI21X1_342
timestamp 1651764895
transform 1 0 984 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_338
timestamp 1651764895
transform -1 0 1096 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_73
timestamp 1651764895
transform 1 0 1096 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_356
timestamp 1651764895
transform -1 0 1192 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_357
timestamp 1651764895
transform -1 0 1256 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_175
timestamp 1651764895
transform 1 0 1256 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_402
timestamp 1651764895
transform 1 0 1320 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_409
timestamp 1651764895
transform -1 0 1432 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_401
timestamp 1651764895
transform -1 0 1480 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_316
timestamp 1651764895
transform 1 0 1480 0 1 4210
box -4 -6 36 206
use INVX1  INVX1_317
timestamp 1651764895
transform -1 0 1544 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_398
timestamp 1651764895
transform 1 0 1544 0 1 4210
box -4 -6 52 206
use FILL  FILL_21_0_0
timestamp 1651764895
transform 1 0 1592 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_1
timestamp 1651764895
transform 1 0 1608 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_0_2
timestamp 1651764895
transform 1 0 1624 0 1 4210
box -4 -6 20 206
use NAND3X1  NAND3X1_408
timestamp 1651764895
transform 1 0 1640 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_400
timestamp 1651764895
transform -1 0 1752 0 1 4210
box -4 -6 52 206
use OAI21X1  OAI21X1_440
timestamp 1651764895
transform 1 0 1752 0 1 4210
box -4 -6 68 206
use AND2X2  AND2X2_74
timestamp 1651764895
transform -1 0 1880 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_345
timestamp 1651764895
transform -1 0 1928 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_361
timestamp 1651764895
transform -1 0 1992 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_183
timestamp 1651764895
transform 1 0 1992 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_362
timestamp 1651764895
transform -1 0 2120 0 1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_35
timestamp 1651764895
transform -1 0 2248 0 1 4210
box -4 -6 132 206
use OAI21X1  OAI21X1_350
timestamp 1651764895
transform 1 0 2248 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_379
timestamp 1651764895
transform 1 0 2312 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_363
timestamp 1651764895
transform -1 0 2440 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_181
timestamp 1651764895
transform 1 0 2440 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_276
timestamp 1651764895
transform 1 0 2504 0 1 4210
box -4 -6 36 206
use AOI21X1  AOI21X1_184
timestamp 1651764895
transform 1 0 2536 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_364
timestamp 1651764895
transform 1 0 2600 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_290
timestamp 1651764895
transform -1 0 2696 0 1 4210
box -4 -6 36 206
use INVX1  INVX1_359
timestamp 1651764895
transform 1 0 2696 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_458
timestamp 1651764895
transform 1 0 2728 0 1 4210
box -4 -6 68 206
use NOR3X1  NOR3X1_46
timestamp 1651764895
transform -1 0 2920 0 1 4210
box -4 -6 132 206
use INVX1  INVX1_323
timestamp 1651764895
transform 1 0 2920 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_429
timestamp 1651764895
transform 1 0 2952 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_508
timestamp 1651764895
transform -1 0 3080 0 1 4210
box -4 -6 68 206
use FILL  FILL_21_1_0
timestamp 1651764895
transform -1 0 3096 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_1
timestamp 1651764895
transform -1 0 3112 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_1_2
timestamp 1651764895
transform -1 0 3128 0 1 4210
box -4 -6 20 206
use NAND3X1  NAND3X1_430
timestamp 1651764895
transform -1 0 3192 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_461
timestamp 1651764895
transform -1 0 3256 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_531
timestamp 1651764895
transform 1 0 3256 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_413
timestamp 1651764895
transform 1 0 3320 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_431
timestamp 1651764895
transform -1 0 3432 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_212
timestamp 1651764895
transform 1 0 3432 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_308
timestamp 1651764895
transform -1 0 3528 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_433
timestamp 1651764895
transform -1 0 3592 0 1 4210
box -4 -6 68 206
use AOI21X1  AOI21X1_220
timestamp 1651764895
transform 1 0 3592 0 1 4210
box -4 -6 68 206
use OAI21X1  OAI21X1_429
timestamp 1651764895
transform 1 0 3656 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_346
timestamp 1651764895
transform 1 0 3720 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_460
timestamp 1651764895
transform 1 0 3752 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_459
timestamp 1651764895
transform 1 0 3816 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_379
timestamp 1651764895
transform 1 0 3880 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_376
timestamp 1651764895
transform 1 0 3928 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_378
timestamp 1651764895
transform 1 0 3976 0 1 4210
box -4 -6 52 206
use NAND3X1  NAND3X1_437
timestamp 1651764895
transform -1 0 4088 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_401
timestamp 1651764895
transform -1 0 4152 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_307
timestamp 1651764895
transform -1 0 4184 0 1 4210
box -4 -6 36 206
use NAND3X1  NAND3X1_534
timestamp 1651764895
transform -1 0 4248 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_538
timestamp 1651764895
transform 1 0 4248 0 1 4210
box -4 -6 52 206
use NAND2X1  NAND2X1_539
timestamp 1651764895
transform -1 0 4344 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_379
timestamp 1651764895
transform -1 0 4376 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_505
timestamp 1651764895
transform -1 0 4440 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_443
timestamp 1651764895
transform -1 0 4488 0 1 4210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_47
timestamp 1651764895
transform -1 0 4600 0 1 4210
box -4 -6 116 206
use INVX1  INVX1_306
timestamp 1651764895
transform 1 0 4600 0 1 4210
box -4 -6 36 206
use FILL  FILL_21_2_0
timestamp 1651764895
transform 1 0 4632 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_1
timestamp 1651764895
transform 1 0 4648 0 1 4210
box -4 -6 20 206
use FILL  FILL_21_2_2
timestamp 1651764895
transform 1 0 4664 0 1 4210
box -4 -6 20 206
use NAND2X1  NAND2X1_368
timestamp 1651764895
transform 1 0 4680 0 1 4210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_42
timestamp 1651764895
transform 1 0 4728 0 1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_366
timestamp 1651764895
transform -1 0 4888 0 1 4210
box -4 -6 52 206
use OR2X2  OR2X2_36
timestamp 1651764895
transform -1 0 4952 0 1 4210
box -4 -6 68 206
use NAND2X1  NAND2X1_365
timestamp 1651764895
transform -1 0 5000 0 1 4210
box -4 -6 52 206
use AND2X2  AND2X2_81
timestamp 1651764895
transform 1 0 5000 0 1 4210
box -4 -6 68 206
use NAND3X1  NAND3X1_384
timestamp 1651764895
transform -1 0 5128 0 1 4210
box -4 -6 68 206
use XOR2X1  XOR2X1_24
timestamp 1651764895
transform 1 0 5128 0 1 4210
box -4 -6 116 206
use NAND2X1  NAND2X1_380
timestamp 1651764895
transform -1 0 5288 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_364
timestamp 1651764895
transform -1 0 5320 0 1 4210
box -4 -6 36 206
use XNOR2X1  XNOR2X1_57
timestamp 1651764895
transform 1 0 5320 0 1 4210
box -4 -6 116 206
use INVX1  INVX1_300
timestamp 1651764895
transform -1 0 5464 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_369
timestamp 1651764895
transform -1 0 5528 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_263
timestamp 1651764895
transform -1 0 5560 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_308
timestamp 1651764895
transform 1 0 5560 0 1 4210
box -4 -6 52 206
use AOI22X1  AOI22X1_43
timestamp 1651764895
transform -1 0 5688 0 1 4210
box -4 -6 84 206
use NAND2X1  NAND2X1_309
timestamp 1651764895
transform 1 0 5688 0 1 4210
box -4 -6 52 206
use XNOR2X1  XNOR2X1_36
timestamp 1651764895
transform 1 0 5736 0 1 4210
box -4 -6 116 206
use INVX1  INVX1_262
timestamp 1651764895
transform 1 0 5848 0 1 4210
box -4 -6 36 206
use NOR2X1  NOR2X1_128
timestamp 1651764895
transform -1 0 5928 0 1 4210
box -4 -6 52 206
use INVX1  INVX1_251
timestamp 1651764895
transform -1 0 5960 0 1 4210
box -4 -6 36 206
use OAI21X1  OAI21X1_357
timestamp 1651764895
transform -1 0 6024 0 1 4210
box -4 -6 68 206
use INVX1  INVX1_250
timestamp 1651764895
transform -1 0 6056 0 1 4210
box -4 -6 36 206
use NAND2X1  NAND2X1_300
timestamp 1651764895
transform -1 0 6104 0 1 4210
box -4 -6 52 206
use NOR2X1  NOR2X1_127
timestamp 1651764895
transform 1 0 6104 0 1 4210
box -4 -6 52 206
use XOR2X1  XOR2X1_40
timestamp 1651764895
transform 1 0 6152 0 1 4210
box -4 -6 116 206
use XNOR2X1  XNOR2X1_62
timestamp 1651764895
transform 1 0 8 0 -1 4610
box -4 -6 116 206
use OAI21X1  OAI21X1_488
timestamp 1651764895
transform 1 0 120 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_509
timestamp 1651764895
transform 1 0 184 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_508
timestamp 1651764895
transform 1 0 232 0 -1 4610
box -4 -6 52 206
use XOR2X1  XOR2X1_29
timestamp 1651764895
transform -1 0 392 0 -1 4610
box -4 -6 116 206
use OAI21X1  OAI21X1_446
timestamp 1651764895
transform 1 0 392 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_464
timestamp 1651764895
transform 1 0 456 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_411
timestamp 1651764895
transform -1 0 584 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_202
timestamp 1651764895
transform 1 0 584 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_484
timestamp 1651764895
transform -1 0 712 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_404
timestamp 1651764895
transform -1 0 760 0 -1 4610
box -4 -6 52 206
use XOR2X1  XOR2X1_30
timestamp 1651764895
transform -1 0 872 0 -1 4610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_44
timestamp 1651764895
transform -1 0 984 0 -1 4610
box -4 -6 116 206
use AOI21X1  AOI21X1_201
timestamp 1651764895
transform 1 0 984 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_413
timestamp 1651764895
transform 1 0 1048 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_200
timestamp 1651764895
transform -1 0 1176 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_174
timestamp 1651764895
transform 1 0 1176 0 -1 4610
box -4 -6 68 206
use NOR3X1  NOR3X1_30
timestamp 1651764895
transform -1 0 1368 0 -1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_344
timestamp 1651764895
transform 1 0 1368 0 -1 4610
box -4 -6 68 206
use AND2X2  AND2X2_91
timestamp 1651764895
transform -1 0 1496 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_403
timestamp 1651764895
transform -1 0 1544 0 -1 4610
box -4 -6 52 206
use FILL  FILL_22_0_0
timestamp 1651764895
transform -1 0 1560 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_1
timestamp 1651764895
transform -1 0 1576 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_0_2
timestamp 1651764895
transform -1 0 1592 0 -1 4610
box -4 -6 20 206
use AOI21X1  AOI21X1_204
timestamp 1651764895
transform -1 0 1656 0 -1 4610
box -4 -6 68 206
use NOR3X1  NOR3X1_31
timestamp 1651764895
transform -1 0 1784 0 -1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_345
timestamp 1651764895
transform 1 0 1784 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_389
timestamp 1651764895
transform 1 0 1848 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_177
timestamp 1651764895
transform 1 0 1912 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_358
timestamp 1651764895
transform 1 0 1976 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_359
timestamp 1651764895
transform -1 0 2104 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_178
timestamp 1651764895
transform 1 0 2104 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_346
timestamp 1651764895
transform 1 0 2168 0 -1 4610
box -4 -6 68 206
use NOR3X1  NOR3X1_32
timestamp 1651764895
transform 1 0 2232 0 -1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_347
timestamp 1651764895
transform -1 0 2424 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_380
timestamp 1651764895
transform 1 0 2424 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_180
timestamp 1651764895
transform -1 0 2552 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_360
timestamp 1651764895
transform 1 0 2552 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_207
timestamp 1651764895
transform -1 0 2680 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_210
timestamp 1651764895
transform -1 0 2744 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_409
timestamp 1651764895
transform 1 0 2744 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_426
timestamp 1651764895
transform 1 0 2792 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_226
timestamp 1651764895
transform 1 0 2856 0 -1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_227
timestamp 1651764895
transform -1 0 2984 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_478
timestamp 1651764895
transform 1 0 2984 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_480
timestamp 1651764895
transform 1 0 3048 0 -1 4610
box -4 -6 52 206
use FILL  FILL_22_1_0
timestamp 1651764895
transform 1 0 3096 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_1
timestamp 1651764895
transform 1 0 3112 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_1_2
timestamp 1651764895
transform 1 0 3128 0 -1 4610
box -4 -6 20 206
use NAND2X1  NAND2X1_482
timestamp 1651764895
transform 1 0 3144 0 -1 4610
box -4 -6 52 206
use AOI21X1  AOI21X1_252
timestamp 1651764895
transform -1 0 3256 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_529
timestamp 1651764895
transform 1 0 3256 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_481
timestamp 1651764895
transform 1 0 3320 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_482
timestamp 1651764895
transform -1 0 3432 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_484
timestamp 1651764895
transform -1 0 3480 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_480
timestamp 1651764895
transform 1 0 3480 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_483
timestamp 1651764895
transform -1 0 3592 0 -1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_484
timestamp 1651764895
transform 1 0 3592 0 -1 4610
box -4 -6 68 206
use NOR3X1  NOR3X1_42
timestamp 1651764895
transform -1 0 3784 0 -1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_408
timestamp 1651764895
transform 1 0 3784 0 -1 4610
box -4 -6 68 206
use INVX1  INVX1_326
timestamp 1651764895
transform -1 0 3880 0 -1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_478
timestamp 1651764895
transform 1 0 3880 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_451
timestamp 1651764895
transform -1 0 3992 0 -1 4610
box -4 -6 52 206
use NOR2X1  NOR2X1_170
timestamp 1651764895
transform -1 0 4040 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_377
timestamp 1651764895
transform 1 0 4040 0 -1 4610
box -4 -6 52 206
use AOI21X1  AOI21X1_216
timestamp 1651764895
transform -1 0 4152 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_436
timestamp 1651764895
transform 1 0 4152 0 -1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_400
timestamp 1651764895
transform 1 0 4216 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_416
timestamp 1651764895
transform -1 0 4328 0 -1 4610
box -4 -6 52 206
use AOI22X1  AOI22X1_46
timestamp 1651764895
transform 1 0 4328 0 -1 4610
box -4 -6 84 206
use INVX1  INVX1_340
timestamp 1651764895
transform 1 0 4408 0 -1 4610
box -4 -6 36 206
use AOI21X1  AOI21X1_217
timestamp 1651764895
transform -1 0 4504 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_373
timestamp 1651764895
transform -1 0 4552 0 -1 4610
box -4 -6 52 206
use AND2X2  AND2X2_92
timestamp 1651764895
transform 1 0 4552 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_370
timestamp 1651764895
transform -1 0 4664 0 -1 4610
box -4 -6 52 206
use FILL  FILL_22_2_0
timestamp 1651764895
transform 1 0 4664 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_1
timestamp 1651764895
transform 1 0 4680 0 -1 4610
box -4 -6 20 206
use FILL  FILL_22_2_2
timestamp 1651764895
transform 1 0 4696 0 -1 4610
box -4 -6 20 206
use NAND2X1  NAND2X1_418
timestamp 1651764895
transform 1 0 4712 0 -1 4610
box -4 -6 52 206
use OAI21X1  OAI21X1_418
timestamp 1651764895
transform -1 0 4824 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_419
timestamp 1651764895
transform -1 0 4872 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_371
timestamp 1651764895
transform -1 0 4920 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_372
timestamp 1651764895
transform -1 0 4968 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_367
timestamp 1651764895
transform -1 0 5016 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_303
timestamp 1651764895
transform 1 0 5016 0 -1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_431
timestamp 1651764895
transform -1 0 5096 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_332
timestamp 1651764895
transform -1 0 5128 0 -1 4610
box -4 -6 36 206
use XOR2X1  XOR2X1_33
timestamp 1651764895
transform -1 0 5240 0 -1 4610
box -4 -6 116 206
use NAND2X1  NAND2X1_361
timestamp 1651764895
transform 1 0 5240 0 -1 4610
box -4 -6 52 206
use AND2X2  AND2X2_93
timestamp 1651764895
transform 1 0 5288 0 -1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_468
timestamp 1651764895
transform -1 0 5416 0 -1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_155
timestamp 1651764895
transform -1 0 5464 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_301
timestamp 1651764895
transform 1 0 5464 0 -1 4610
box -4 -6 36 206
use AND2X2  AND2X2_83
timestamp 1651764895
transform 1 0 5496 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_421
timestamp 1651764895
transform 1 0 5560 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_360
timestamp 1651764895
transform -1 0 5656 0 -1 4610
box -4 -6 52 206
use INVX1  INVX1_302
timestamp 1651764895
transform -1 0 5688 0 -1 4610
box -4 -6 36 206
use AND2X2  AND2X2_94
timestamp 1651764895
transform -1 0 5752 0 -1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_358
timestamp 1651764895
transform 1 0 5752 0 -1 4610
box -4 -6 52 206
use AOI22X1  AOI22X1_52
timestamp 1651764895
transform -1 0 5880 0 -1 4610
box -4 -6 84 206
use NAND2X1  NAND2X1_307
timestamp 1651764895
transform -1 0 5928 0 -1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_357
timestamp 1651764895
transform -1 0 5976 0 -1 4610
box -4 -6 52 206
use AND2X2  AND2X2_95
timestamp 1651764895
transform 1 0 5976 0 -1 4610
box -4 -6 68 206
use NOR3X1  NOR3X1_43
timestamp 1651764895
transform 1 0 6040 0 -1 4610
box -4 -6 132 206
use NAND2X1  NAND2X1_304
timestamp 1651764895
transform -1 0 6216 0 -1 4610
box -4 -6 52 206
use FILL  FILL_23_1
timestamp 1651764895
transform -1 0 6232 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_2
timestamp 1651764895
transform -1 0 6248 0 -1 4610
box -4 -6 20 206
use FILL  FILL_23_3
timestamp 1651764895
transform -1 0 6264 0 -1 4610
box -4 -6 20 206
use XOR2X1  XOR2X1_49
timestamp 1651764895
transform 1 0 8 0 1 4610
box -4 -6 116 206
use AND2X2  AND2X2_106
timestamp 1651764895
transform -1 0 184 0 1 4610
box -4 -6 68 206
use NOR2X1  NOR2X1_187
timestamp 1651764895
transform -1 0 232 0 1 4610
box -4 -6 52 206
use XOR2X1  XOR2X1_46
timestamp 1651764895
transform -1 0 344 0 1 4610
box -4 -6 116 206
use XNOR2X1  XNOR2X1_68
timestamp 1651764895
transform -1 0 456 0 1 4610
box -4 -6 116 206
use NAND3X1  NAND3X1_512
timestamp 1651764895
transform -1 0 520 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_464
timestamp 1651764895
transform -1 0 568 0 1 4610
box -4 -6 52 206
use XNOR2X1  XNOR2X1_50
timestamp 1651764895
transform -1 0 680 0 1 4610
box -4 -6 116 206
use XOR2X1  XOR2X1_36
timestamp 1651764895
transform 1 0 680 0 1 4610
box -4 -6 116 206
use NOR3X1  NOR3X1_36
timestamp 1651764895
transform -1 0 920 0 1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_398
timestamp 1651764895
transform 1 0 920 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_320
timestamp 1651764895
transform -1 0 1016 0 1 4610
box -4 -6 36 206
use INVX1  INVX1_29
timestamp 1651764895
transform 1 0 1016 0 1 4610
box -4 -6 36 206
use NOR2X1  NOR2X1_175
timestamp 1651764895
transform 1 0 1048 0 1 4610
box -4 -6 52 206
use NOR3X1  NOR3X1_37
timestamp 1651764895
transform -1 0 1224 0 1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_400
timestamp 1651764895
transform 1 0 1224 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_321
timestamp 1651764895
transform 1 0 1288 0 1 4610
box -4 -6 36 206
use AOI21X1  AOI21X1_203
timestamp 1651764895
transform 1 0 1320 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_414
timestamp 1651764895
transform 1 0 1384 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_205
timestamp 1651764895
transform 1 0 1448 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_415
timestamp 1651764895
transform 1 0 1512 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_0_0
timestamp 1651764895
transform 1 0 1576 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_1
timestamp 1651764895
transform 1 0 1592 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_0_2
timestamp 1651764895
transform 1 0 1608 0 1 4610
box -4 -6 20 206
use NOR3X1  NOR3X1_38
timestamp 1651764895
transform 1 0 1624 0 1 4610
box -4 -6 132 206
use OAI21X1  OAI21X1_399
timestamp 1651764895
transform 1 0 1752 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_416
timestamp 1651764895
transform -1 0 1880 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_206
timestamp 1651764895
transform 1 0 1880 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_347
timestamp 1651764895
transform -1 0 2008 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_349
timestamp 1651764895
transform 1 0 2008 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_242
timestamp 1651764895
transform 1 0 2072 0 1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_348
timestamp 1651764895
transform -1 0 2168 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_336
timestamp 1651764895
transform 1 0 2168 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_283
timestamp 1651764895
transform 1 0 2216 0 1 4610
box -4 -6 52 206
use NOR3X1  NOR3X1_33
timestamp 1651764895
transform -1 0 2392 0 1 4610
box -4 -6 132 206
use INVX1  INVX1_282
timestamp 1651764895
transform 1 0 2392 0 1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_425
timestamp 1651764895
transform -1 0 2488 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_422
timestamp 1651764895
transform -1 0 2552 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_420
timestamp 1651764895
transform 1 0 2552 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_424
timestamp 1651764895
transform -1 0 2680 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_423
timestamp 1651764895
transform -1 0 2744 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_253
timestamp 1651764895
transform 1 0 2744 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_479
timestamp 1651764895
transform 1 0 2808 0 1 4610
box -4 -6 52 206
use NOR3X1  NOR3X1_45
timestamp 1651764895
transform -1 0 2984 0 1 4610
box -4 -6 132 206
use NAND3X1  NAND3X1_481
timestamp 1651764895
transform 1 0 2984 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_503
timestamp 1651764895
transform -1 0 3112 0 1 4610
box -4 -6 68 206
use FILL  FILL_23_1_0
timestamp 1651764895
transform -1 0 3128 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_1
timestamp 1651764895
transform -1 0 3144 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_1_2
timestamp 1651764895
transform -1 0 3160 0 1 4610
box -4 -6 20 206
use INVX1  INVX1_377
timestamp 1651764895
transform -1 0 3192 0 1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_485
timestamp 1651764895
transform -1 0 3256 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_229
timestamp 1651764895
transform 1 0 3256 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_348
timestamp 1651764895
transform 1 0 3320 0 1 4610
box -4 -6 36 206
use AOI21X1  AOI21X1_230
timestamp 1651764895
transform -1 0 3416 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_483
timestamp 1651764895
transform 1 0 3416 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_460
timestamp 1651764895
transform 1 0 3480 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_461
timestamp 1651764895
transform 1 0 3544 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_434
timestamp 1651764895
transform -1 0 3672 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_213
timestamp 1651764895
transform 1 0 3672 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_438
timestamp 1651764895
transform -1 0 3800 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_435
timestamp 1651764895
transform -1 0 3864 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_327
timestamp 1651764895
transform -1 0 3896 0 1 4610
box -4 -6 36 206
use OAI21X1  OAI21X1_409
timestamp 1651764895
transform -1 0 3960 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_410
timestamp 1651764895
transform 1 0 3960 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_439
timestamp 1651764895
transform -1 0 4088 0 1 4610
box -4 -6 68 206
use AOI22X1  AOI22X1_47
timestamp 1651764895
transform -1 0 4168 0 1 4610
box -4 -6 84 206
use NAND2X1  NAND2X1_417
timestamp 1651764895
transform 1 0 4168 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_440
timestamp 1651764895
transform -1 0 4280 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_443
timestamp 1651764895
transform -1 0 4344 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_441
timestamp 1651764895
transform -1 0 4408 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_411
timestamp 1651764895
transform 1 0 4408 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_412
timestamp 1651764895
transform 1 0 4472 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_442
timestamp 1651764895
transform -1 0 4600 0 1 4610
box -4 -6 68 206
use AOI22X1  AOI22X1_49
timestamp 1651764895
transform -1 0 4680 0 1 4610
box -4 -6 84 206
use FILL  FILL_23_2_0
timestamp 1651764895
transform 1 0 4680 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_1
timestamp 1651764895
transform 1 0 4696 0 1 4610
box -4 -6 20 206
use FILL  FILL_23_2_2
timestamp 1651764895
transform 1 0 4712 0 1 4610
box -4 -6 20 206
use NAND2X1  NAND2X1_420
timestamp 1651764895
transform 1 0 4728 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_444
timestamp 1651764895
transform 1 0 4776 0 1 4610
box -4 -6 68 206
use AOI22X1  AOI22X1_48
timestamp 1651764895
transform -1 0 4920 0 1 4610
box -4 -6 84 206
use INVX1  INVX1_331
timestamp 1651764895
transform 1 0 4920 0 1 4610
box -4 -6 36 206
use NAND2X1  NAND2X1_432
timestamp 1651764895
transform -1 0 5000 0 1 4610
box -4 -6 52 206
use NAND2X1  NAND2X1_433
timestamp 1651764895
transform -1 0 5048 0 1 4610
box -4 -6 52 206
use NAND3X1  NAND3X1_495
timestamp 1651764895
transform -1 0 5112 0 1 4610
box -4 -6 68 206
use XNOR2X1  XNOR2X1_46
timestamp 1651764895
transform -1 0 5224 0 1 4610
box -4 -6 116 206
use OAI21X1  OAI21X1_414
timestamp 1651764895
transform 1 0 5224 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_413
timestamp 1651764895
transform 1 0 5288 0 1 4610
box -4 -6 68 206
use OR2X2  OR2X2_41
timestamp 1651764895
transform 1 0 5352 0 1 4610
box -4 -6 68 206
use NAND2X1  NAND2X1_422
timestamp 1651764895
transform -1 0 5464 0 1 4610
box -4 -6 52 206
use AOI22X1  AOI22X1_51
timestamp 1651764895
transform 1 0 5464 0 1 4610
box -4 -6 84 206
use AOI22X1  AOI22X1_50
timestamp 1651764895
transform -1 0 5624 0 1 4610
box -4 -6 84 206
use OR2X2  OR2X2_35
timestamp 1651764895
transform -1 0 5688 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_416
timestamp 1651764895
transform 1 0 5688 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_415
timestamp 1651764895
transform 1 0 5752 0 1 4610
box -4 -6 68 206
use NAND3X1  NAND3X1_452
timestamp 1651764895
transform -1 0 5880 0 1 4610
box -4 -6 68 206
use INVX1  INVX1_329
timestamp 1651764895
transform -1 0 5912 0 1 4610
box -4 -6 36 206
use NAND3X1  NAND3X1_450
timestamp 1651764895
transform 1 0 5912 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_308
timestamp 1651764895
transform -1 0 6040 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_214
timestamp 1651764895
transform 1 0 6040 0 1 4610
box -4 -6 68 206
use OAI21X1  OAI21X1_417
timestamp 1651764895
transform -1 0 6168 0 1 4610
box -4 -6 68 206
use AOI21X1  AOI21X1_215
timestamp 1651764895
transform -1 0 6232 0 1 4610
box -4 -6 68 206
use FILL  FILL_24_1
timestamp 1651764895
transform 1 0 6232 0 1 4610
box -4 -6 20 206
use FILL  FILL_24_2
timestamp 1651764895
transform 1 0 6248 0 1 4610
box -4 -6 20 206
use XNOR2X1  XNOR2X1_75
timestamp 1651764895
transform 1 0 8 0 -1 5010
box -4 -6 116 206
use NAND2X1  NAND2X1_520
timestamp 1651764895
transform -1 0 168 0 -1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_193
timestamp 1651764895
transform -1 0 216 0 -1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_74
timestamp 1651764895
transform -1 0 328 0 -1 5010
box -4 -6 116 206
use NAND2X1  NAND2X1_515
timestamp 1651764895
transform -1 0 376 0 -1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_190
timestamp 1651764895
transform -1 0 424 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_372
timestamp 1651764895
transform 1 0 424 0 -1 5010
box -4 -6 36 206
use AND2X2  AND2X2_105
timestamp 1651764895
transform -1 0 520 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_506
timestamp 1651764895
transform 1 0 520 0 -1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_65
timestamp 1651764895
transform -1 0 680 0 -1 5010
box -4 -6 116 206
use NAND2X1  NAND2X1_505
timestamp 1651764895
transform -1 0 728 0 -1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_64
timestamp 1651764895
transform 1 0 728 0 -1 5010
box -4 -6 116 206
use NAND2X1  NAND2X1_503
timestamp 1651764895
transform 1 0 840 0 -1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_387
timestamp 1651764895
transform -1 0 936 0 -1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_457
timestamp 1651764895
transform -1 0 984 0 -1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_220
timestamp 1651764895
transform 1 0 984 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_174
timestamp 1651764895
transform 1 0 1032 0 -1 5010
box -4 -6 36 206
use INVX1  INVX1_203
timestamp 1651764895
transform 1 0 1064 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_221
timestamp 1651764895
transform 1 0 1096 0 -1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_102
timestamp 1651764895
transform 1 0 1160 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_204
timestamp 1651764895
transform 1 0 1208 0 -1 5010
box -4 -6 36 206
use AND2X2  AND2X2_49
timestamp 1651764895
transform 1 0 1240 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_270
timestamp 1651764895
transform 1 0 1304 0 -1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_119
timestamp 1651764895
transform 1 0 1368 0 -1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_441
timestamp 1651764895
transform -1 0 1480 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_401
timestamp 1651764895
transform 1 0 1480 0 -1 5010
box -4 -6 68 206
use FILL  FILL_24_0_0
timestamp 1651764895
transform 1 0 1544 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_1
timestamp 1651764895
transform 1 0 1560 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_0_2
timestamp 1651764895
transform 1 0 1576 0 -1 5010
box -4 -6 20 206
use NOR3X1  NOR3X1_39
timestamp 1651764895
transform 1 0 1592 0 -1 5010
box -4 -6 132 206
use XOR2X1  XOR2X1_38
timestamp 1651764895
transform 1 0 1720 0 -1 5010
box -4 -6 116 206
use INVX1  INVX1_280
timestamp 1651764895
transform 1 0 1832 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_330
timestamp 1651764895
transform 1 0 1864 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_279
timestamp 1651764895
transform 1 0 1928 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_329
timestamp 1651764895
transform 1 0 1960 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_350
timestamp 1651764895
transform -1 0 2088 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_382
timestamp 1651764895
transform 1 0 2088 0 -1 5010
box -4 -6 52 206
use AOI21X1  AOI21X1_208
timestamp 1651764895
transform 1 0 2136 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_417
timestamp 1651764895
transform -1 0 2264 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_418
timestamp 1651764895
transform -1 0 2328 0 -1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_209
timestamp 1651764895
transform 1 0 2328 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_419
timestamp 1651764895
transform -1 0 2456 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_421
timestamp 1651764895
transform -1 0 2520 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_405
timestamp 1651764895
transform -1 0 2584 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_404
timestamp 1651764895
transform -1 0 2648 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_430
timestamp 1651764895
transform 1 0 2648 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_454
timestamp 1651764895
transform -1 0 2776 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_456
timestamp 1651764895
transform 1 0 2776 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_358
timestamp 1651764895
transform -1 0 2872 0 -1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_457
timestamp 1651764895
transform -1 0 2936 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_455
timestamp 1651764895
transform -1 0 3000 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_478
timestamp 1651764895
transform 1 0 3000 0 -1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_61
timestamp 1651764895
transform 1 0 3048 0 -1 5010
box -4 -6 116 206
use FILL  FILL_24_1_0
timestamp 1651764895
transform 1 0 3160 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_1
timestamp 1651764895
transform 1 0 3176 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_1_2
timestamp 1651764895
transform 1 0 3192 0 -1 5010
box -4 -6 20 206
use NAND3X1  NAND3X1_528
timestamp 1651764895
transform 1 0 3208 0 -1 5010
box -4 -6 68 206
use XOR2X1  XOR2X1_43
timestamp 1651764895
transform 1 0 3272 0 -1 5010
box -4 -6 116 206
use NAND3X1  NAND3X1_507
timestamp 1651764895
transform -1 0 3448 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_480
timestamp 1651764895
transform 1 0 3448 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_509
timestamp 1651764895
transform 1 0 3512 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_370
timestamp 1651764895
transform 1 0 3576 0 -1 5010
box -4 -6 36 206
use INVX1  INVX1_362
timestamp 1651764895
transform 1 0 3608 0 -1 5010
box -4 -6 36 206
use NAND3X1  NAND3X1_487
timestamp 1651764895
transform 1 0 3640 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_486
timestamp 1651764895
transform 1 0 3704 0 -1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_231
timestamp 1651764895
transform 1 0 3768 0 -1 5010
box -4 -6 68 206
use AOI22X1  AOI22X1_55
timestamp 1651764895
transform -1 0 3912 0 -1 5010
box -4 -6 84 206
use NAND2X1  NAND2X1_453
timestamp 1651764895
transform -1 0 3960 0 -1 5010
box -4 -6 52 206
use AOI22X1  AOI22X1_54
timestamp 1651764895
transform -1 0 4040 0 -1 5010
box -4 -6 84 206
use OAI21X1  OAI21X1_464
timestamp 1651764895
transform -1 0 4104 0 -1 5010
box -4 -6 68 206
use AND2X2  AND2X2_109
timestamp 1651764895
transform -1 0 4168 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_540
timestamp 1651764895
transform -1 0 4216 0 -1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_465
timestamp 1651764895
transform 1 0 4216 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_341
timestamp 1651764895
transform -1 0 4312 0 -1 5010
box -4 -6 36 206
use AOI21X1  AOI21X1_233
timestamp 1651764895
transform 1 0 4312 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_489
timestamp 1651764895
transform -1 0 4440 0 -1 5010
box -4 -6 68 206
use OR2X2  OR2X2_47
timestamp 1651764895
transform 1 0 4440 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_456
timestamp 1651764895
transform -1 0 4568 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_445
timestamp 1651764895
transform 1 0 4568 0 -1 5010
box -4 -6 52 206
use INVX1  INVX1_339
timestamp 1651764895
transform -1 0 4648 0 -1 5010
box -4 -6 36 206
use FILL  FILL_24_2_0
timestamp 1651764895
transform -1 0 4664 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_1
timestamp 1651764895
transform -1 0 4680 0 -1 5010
box -4 -6 20 206
use FILL  FILL_24_2_2
timestamp 1651764895
transform -1 0 4696 0 -1 5010
box -4 -6 20 206
use NAND2X1  NAND2X1_444
timestamp 1651764895
transform -1 0 4744 0 -1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_171
timestamp 1651764895
transform 1 0 4744 0 -1 5010
box -4 -6 52 206
use AND2X2  AND2X2_99
timestamp 1651764895
transform 1 0 4792 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_425
timestamp 1651764895
transform 1 0 4856 0 -1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_241
timestamp 1651764895
transform -1 0 4984 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_434
timestamp 1651764895
transform -1 0 5032 0 -1 5010
box -4 -6 52 206
use AND2X2  AND2X2_102
timestamp 1651764895
transform 1 0 5032 0 -1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_473
timestamp 1651764895
transform 1 0 5096 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_486
timestamp 1651764895
transform 1 0 5160 0 -1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_493
timestamp 1651764895
transform -1 0 5256 0 -1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_477
timestamp 1651764895
transform -1 0 5320 0 -1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_180
timestamp 1651764895
transform -1 0 5368 0 -1 5010
box -4 -6 52 206
use NAND3X1  NAND3X1_445
timestamp 1651764895
transform 1 0 5368 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_446
timestamp 1651764895
transform 1 0 5432 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_424
timestamp 1651764895
transform 1 0 5496 0 -1 5010
box -4 -6 52 206
use NAND3X1  NAND3X1_448
timestamp 1651764895
transform -1 0 5608 0 -1 5010
box -4 -6 68 206
use INVX1  INVX1_328
timestamp 1651764895
transform 1 0 5608 0 -1 5010
box -4 -6 36 206
use NAND3X1  NAND3X1_447
timestamp 1651764895
transform 1 0 5640 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_449
timestamp 1651764895
transform -1 0 5768 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_451
timestamp 1651764895
transform -1 0 5832 0 -1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_239
timestamp 1651764895
transform 1 0 5832 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_453
timestamp 1651764895
transform -1 0 5960 0 -1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_454
timestamp 1651764895
transform 1 0 5960 0 -1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_423
timestamp 1651764895
transform 1 0 6024 0 -1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_60
timestamp 1651764895
transform 1 0 6072 0 -1 5010
box -4 -6 116 206
use NAND3X1  NAND3X1_328
timestamp 1651764895
transform 1 0 6184 0 -1 5010
box -4 -6 68 206
use FILL  FILL_25_1
timestamp 1651764895
transform -1 0 6264 0 -1 5010
box -4 -6 20 206
use NAND2X1  NAND2X1_519
timestamp 1651764895
transform 1 0 8 0 1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_194
timestamp 1651764895
transform -1 0 104 0 1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_73
timestamp 1651764895
transform 1 0 104 0 1 5010
box -4 -6 116 206
use OAI21X1  OAI21X1_493
timestamp 1651764895
transform -1 0 280 0 1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_189
timestamp 1651764895
transform -1 0 328 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_516
timestamp 1651764895
transform -1 0 376 0 1 5010
box -4 -6 52 206
use OAI22X1  OAI22X1_11
timestamp 1651764895
transform 1 0 376 0 1 5010
box -4 -6 84 206
use NOR2X1  NOR2X1_192
timestamp 1651764895
transform -1 0 504 0 1 5010
box -4 -6 52 206
use NOR2X1  NOR2X1_191
timestamp 1651764895
transform -1 0 552 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_504
timestamp 1651764895
transform 1 0 552 0 1 5010
box -4 -6 52 206
use XNOR2X1  XNOR2X1_66
timestamp 1651764895
transform -1 0 712 0 1 5010
box -4 -6 116 206
use NAND2X1  NAND2X1_458
timestamp 1651764895
transform -1 0 760 0 1 5010
box -4 -6 52 206
use OR2X2  OR2X2_49
timestamp 1651764895
transform 1 0 760 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_486
timestamp 1651764895
transform -1 0 888 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_459
timestamp 1651764895
transform -1 0 936 0 1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_438
timestamp 1651764895
transform 1 0 936 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_439
timestamp 1651764895
transform -1 0 1064 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_437
timestamp 1651764895
transform -1 0 1128 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_383
timestamp 1651764895
transform -1 0 1192 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_388
timestamp 1651764895
transform -1 0 1240 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_219
timestamp 1651764895
transform -1 0 1288 0 1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_268
timestamp 1651764895
transform 1 0 1288 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_324
timestamp 1651764895
transform 1 0 1352 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_269
timestamp 1651764895
transform 1 0 1416 0 1 5010
box -4 -6 68 206
use XOR2X1  XOR2X1_17
timestamp 1651764895
transform 1 0 1480 0 1 5010
box -4 -6 116 206
use FILL  FILL_25_0_0
timestamp 1651764895
transform 1 0 1592 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_0_1
timestamp 1651764895
transform 1 0 1608 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_0_2
timestamp 1651764895
transform 1 0 1624 0 1 5010
box -4 -6 20 206
use NOR2X1  NOR2X1_140
timestamp 1651764895
transform 1 0 1640 0 1 5010
box -4 -6 52 206
use AOI21X1  AOI21X1_164
timestamp 1651764895
transform -1 0 1752 0 1 5010
box -4 -6 68 206
use NOR2X1  NOR2X1_118
timestamp 1651764895
transform -1 0 1800 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_472
timestamp 1651764895
transform 1 0 1800 0 1 5010
box -4 -6 52 206
use OR2X2  OR2X2_53
timestamp 1651764895
transform 1 0 1848 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_473
timestamp 1651764895
transform 1 0 1912 0 1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_483
timestamp 1651764895
transform -1 0 2024 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_353
timestamp 1651764895
transform -1 0 2056 0 1 5010
box -4 -6 36 206
use NAND2X1  NAND2X1_476
timestamp 1651764895
transform -1 0 2104 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_471
timestamp 1651764895
transform 1 0 2104 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_475
timestamp 1651764895
transform -1 0 2200 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_474
timestamp 1651764895
transform -1 0 2248 0 1 5010
box -4 -6 52 206
use INVX1  INVX1_315
timestamp 1651764895
transform -1 0 2280 0 1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_402
timestamp 1651764895
transform -1 0 2344 0 1 5010
box -4 -6 68 206
use NOR3X1  NOR3X1_40
timestamp 1651764895
transform -1 0 2472 0 1 5010
box -4 -6 132 206
use OAI21X1  OAI21X1_431
timestamp 1651764895
transform 1 0 2472 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_322
timestamp 1651764895
transform 1 0 2536 0 1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_403
timestamp 1651764895
transform 1 0 2568 0 1 5010
box -4 -6 68 206
use NOR3X1  NOR3X1_41
timestamp 1651764895
transform 1 0 2632 0 1 5010
box -4 -6 132 206
use AOI21X1  AOI21X1_222
timestamp 1651764895
transform -1 0 2824 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_224
timestamp 1651764895
transform 1 0 2824 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_357
timestamp 1651764895
transform -1 0 2920 0 1 5010
box -4 -6 36 206
use AOI21X1  AOI21X1_223
timestamp 1651764895
transform -1 0 2984 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_225
timestamp 1651764895
transform -1 0 3048 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_529
timestamp 1651764895
transform -1 0 3096 0 1 5010
box -4 -6 52 206
use FILL  FILL_25_1_0
timestamp 1651764895
transform 1 0 3096 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_1_1
timestamp 1651764895
transform 1 0 3112 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_1_2
timestamp 1651764895
transform 1 0 3128 0 1 5010
box -4 -6 20 206
use AND2X2  AND2X2_108
timestamp 1651764895
transform 1 0 3144 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_499
timestamp 1651764895
transform 1 0 3208 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_498
timestamp 1651764895
transform -1 0 3304 0 1 5010
box -4 -6 52 206
use NAND3X1  NAND3X1_510
timestamp 1651764895
transform -1 0 3368 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_497
timestamp 1651764895
transform -1 0 3416 0 1 5010
box -4 -6 52 206
use NAND2X1  NAND2X1_533
timestamp 1651764895
transform 1 0 3416 0 1 5010
box -4 -6 52 206
use NAND3X1  NAND3X1_533
timestamp 1651764895
transform -1 0 3528 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_255
timestamp 1651764895
transform -1 0 3592 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_500
timestamp 1651764895
transform 1 0 3592 0 1 5010
box -4 -6 52 206
use AOI21X1  AOI21X1_256
timestamp 1651764895
transform 1 0 3640 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_532
timestamp 1651764895
transform 1 0 3704 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_232
timestamp 1651764895
transform 1 0 3768 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_506
timestamp 1651764895
transform -1 0 3896 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_369
timestamp 1651764895
transform 1 0 3896 0 1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_479
timestamp 1651764895
transform -1 0 3992 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_463
timestamp 1651764895
transform 1 0 3992 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_347
timestamp 1651764895
transform 1 0 4056 0 1 5010
box -4 -6 36 206
use OAI21X1  OAI21X1_462
timestamp 1651764895
transform 1 0 4088 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_234
timestamp 1651764895
transform 1 0 4152 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_488
timestamp 1651764895
transform 1 0 4216 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_466
timestamp 1651764895
transform 1 0 4280 0 1 5010
box -4 -6 68 206
use OAI21X1  OAI21X1_467
timestamp 1651764895
transform 1 0 4344 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_363
timestamp 1651764895
transform -1 0 4440 0 1 5010
box -4 -6 36 206
use NAND3X1  NAND3X1_492
timestamp 1651764895
transform -1 0 4504 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_490
timestamp 1651764895
transform -1 0 4568 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_258
timestamp 1651764895
transform -1 0 4632 0 1 5010
box -4 -6 68 206
use FILL  FILL_25_2_0
timestamp 1651764895
transform -1 0 4648 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_2_1
timestamp 1651764895
transform -1 0 4664 0 1 5010
box -4 -6 20 206
use FILL  FILL_25_2_2
timestamp 1651764895
transform -1 0 4680 0 1 5010
box -4 -6 20 206
use NAND3X1  NAND3X1_491
timestamp 1651764895
transform -1 0 4744 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_236
timestamp 1651764895
transform 1 0 4744 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_497
timestamp 1651764895
transform 1 0 4808 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_498
timestamp 1651764895
transform 1 0 4872 0 1 5010
box -4 -6 68 206
use AOI21X1  AOI21X1_235
timestamp 1651764895
transform 1 0 4936 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_493
timestamp 1651764895
transform 1 0 5000 0 1 5010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_58
timestamp 1651764895
transform 1 0 5064 0 1 5010
box -4 -6 116 206
use INVX1  INVX1_366
timestamp 1651764895
transform -1 0 5208 0 1 5010
box -4 -6 36 206
use OR2X2  OR2X2_54
timestamp 1651764895
transform -1 0 5272 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_367
timestamp 1651764895
transform -1 0 5304 0 1 5010
box -4 -6 36 206
use XNOR2X1  XNOR2X1_82
timestamp 1651764895
transform -1 0 5416 0 1 5010
box -4 -6 116 206
use NAND3X1  NAND3X1_496
timestamp 1651764895
transform 1 0 5416 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_500
timestamp 1651764895
transform 1 0 5480 0 1 5010
box -4 -6 68 206
use AND2X2  AND2X2_103
timestamp 1651764895
transform -1 0 5608 0 1 5010
box -4 -6 68 206
use INVX1  INVX1_330
timestamp 1651764895
transform -1 0 5640 0 1 5010
box -4 -6 36 206
use NAND3X1  NAND3X1_501
timestamp 1651764895
transform 1 0 5640 0 1 5010
box -4 -6 68 206
use NAND3X1  NAND3X1_504
timestamp 1651764895
transform 1 0 5704 0 1 5010
box -4 -6 68 206
use AND2X2  AND2X2_96
timestamp 1651764895
transform -1 0 5832 0 1 5010
box -4 -6 68 206
use NAND2X1  NAND2X1_487
timestamp 1651764895
transform 1 0 5832 0 1 5010
box -4 -6 52 206
use OAI21X1  OAI21X1_472
timestamp 1651764895
transform 1 0 5880 0 1 5010
box -4 -6 68 206
use XOR2X1  XOR2X1_32
timestamp 1651764895
transform -1 0 6056 0 1 5010
box -4 -6 116 206
use INVX1  INVX1_227
timestamp 1651764895
transform -1 0 6088 0 1 5010
box -4 -6 36 206
use XOR2X1  XOR2X1_42
timestamp 1651764895
transform 1 0 6088 0 1 5010
box -4 -6 116 206
use NAND3X1  NAND3X1_337
timestamp 1651764895
transform 1 0 6200 0 1 5010
box -4 -6 68 206
use AOI22X1  AOI22X1_58
timestamp 1651764895
transform -1 0 88 0 -1 5410
box -4 -6 84 206
use AOI21X1  AOI21X1_244
timestamp 1651764895
transform 1 0 88 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_490
timestamp 1651764895
transform 1 0 152 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_373
timestamp 1651764895
transform 1 0 216 0 -1 5410
box -4 -6 36 206
use AOI21X1  AOI21X1_245
timestamp 1651764895
transform -1 0 312 0 -1 5410
box -4 -6 68 206
use AOI22X1  AOI22X1_57
timestamp 1651764895
transform 1 0 312 0 -1 5410
box -4 -6 84 206
use NAND2X1  NAND2X1_514
timestamp 1651764895
transform -1 0 440 0 -1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_517
timestamp 1651764895
transform -1 0 488 0 -1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_518
timestamp 1651764895
transform -1 0 536 0 -1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_513
timestamp 1651764895
transform 1 0 536 0 -1 5410
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1651764895
transform -1 0 616 0 -1 5410
box -4 -6 36 206
use XNOR2X1  XNOR2X1_76
timestamp 1651764895
transform 1 0 616 0 -1 5410
box -4 -6 116 206
use XOR2X1  XOR2X1_44
timestamp 1651764895
transform -1 0 840 0 -1 5410
box -4 -6 116 206
use AOI21X1  AOI21X1_243
timestamp 1651764895
transform -1 0 904 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_371
timestamp 1651764895
transform -1 0 936 0 -1 5410
box -4 -6 36 206
use XOR2X1  XOR2X1_34
timestamp 1651764895
transform -1 0 1048 0 -1 5410
box -4 -6 116 206
use INVX1  INVX1_241
timestamp 1651764895
transform -1 0 1080 0 -1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_436
timestamp 1651764895
transform -1 0 1144 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_384
timestamp 1651764895
transform -1 0 1208 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_332
timestamp 1651764895
transform 1 0 1208 0 -1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_281
timestamp 1651764895
transform -1 0 1304 0 -1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_334
timestamp 1651764895
transform 1 0 1304 0 -1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_325
timestamp 1651764895
transform 1 0 1352 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_326
timestamp 1651764895
transform 1 0 1416 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_335
timestamp 1651764895
transform -1 0 1528 0 -1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_141
timestamp 1651764895
transform 1 0 1528 0 -1 5410
box -4 -6 52 206
use FILL  FILL_26_0_0
timestamp 1651764895
transform 1 0 1576 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_0_1
timestamp 1651764895
transform 1 0 1592 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_0_2
timestamp 1651764895
transform 1 0 1608 0 -1 5410
box -4 -6 20 206
use NAND3X1  NAND3X1_344
timestamp 1651764895
transform 1 0 1624 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_278
timestamp 1651764895
transform 1 0 1688 0 -1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_345
timestamp 1651764895
transform 1 0 1720 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_346
timestamp 1651764895
transform -1 0 1848 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_165
timestamp 1651764895
transform 1 0 1848 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_383
timestamp 1651764895
transform 1 0 1912 0 -1 5410
box -4 -6 52 206
use INVX1  INVX1_354
timestamp 1651764895
transform 1 0 1960 0 -1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_469
timestamp 1651764895
transform 1 0 1992 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_466
timestamp 1651764895
transform -1 0 2120 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_468
timestamp 1651764895
transform 1 0 2120 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_248
timestamp 1651764895
transform 1 0 2184 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_465
timestamp 1651764895
transform 1 0 2248 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_221
timestamp 1651764895
transform 1 0 2312 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_470
timestamp 1651764895
transform 1 0 2376 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_527
timestamp 1651764895
transform 1 0 2440 0 -1 5410
box -4 -6 52 206
use NOR3X1  NOR3X1_44
timestamp 1651764895
transform -1 0 2616 0 -1 5410
box -4 -6 132 206
use OAI21X1  OAI21X1_453
timestamp 1651764895
transform 1 0 2616 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_476
timestamp 1651764895
transform 1 0 2680 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_474
timestamp 1651764895
transform -1 0 2808 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_249
timestamp 1651764895
transform -1 0 2872 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_472
timestamp 1651764895
transform 1 0 2872 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_475
timestamp 1651764895
transform 1 0 2936 0 -1 5410
box -4 -6 68 206
use AND2X2  AND2X2_107
timestamp 1651764895
transform 1 0 3000 0 -1 5410
box -4 -6 68 206
use NOR2X1  NOR2X1_195
timestamp 1651764895
transform -1 0 3112 0 -1 5410
box -4 -6 52 206
use FILL  FILL_26_1_0
timestamp 1651764895
transform -1 0 3128 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_1_1
timestamp 1651764895
transform -1 0 3144 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_1_2
timestamp 1651764895
transform -1 0 3160 0 -1 5410
box -4 -6 20 206
use OAI22X1  OAI22X1_13
timestamp 1651764895
transform -1 0 3240 0 -1 5410
box -4 -6 84 206
use NAND3X1  NAND3X1_524
timestamp 1651764895
transform -1 0 3304 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_528
timestamp 1651764895
transform -1 0 3352 0 -1 5410
box -4 -6 52 206
use OR2X2  OR2X2_58
timestamp 1651764895
transform 1 0 3352 0 -1 5410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_59
timestamp 1651764895
transform 1 0 3416 0 -1 5410
box -4 -6 116 206
use XOR2X1  XOR2X1_52
timestamp 1651764895
transform -1 0 3640 0 -1 5410
box -4 -6 116 206
use NAND2X1  NAND2X1_496
timestamp 1651764895
transform 1 0 3640 0 -1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_507
timestamp 1651764895
transform 1 0 3688 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_257
timestamp 1651764895
transform 1 0 3752 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_535
timestamp 1651764895
transform 1 0 3816 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_508
timestamp 1651764895
transform 1 0 3880 0 -1 5410
box -4 -6 68 206
use NOR3X1  NOR3X1_49
timestamp 1651764895
transform 1 0 3944 0 -1 5410
box -4 -6 132 206
use NAND3X1  NAND3X1_536
timestamp 1651764895
transform -1 0 4136 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_260
timestamp 1651764895
transform 1 0 4136 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_512
timestamp 1651764895
transform 1 0 4200 0 -1 5410
box -4 -6 68 206
use NOR3X1  NOR3X1_50
timestamp 1651764895
transform 1 0 4264 0 -1 5410
box -4 -6 132 206
use AOI21X1  AOI21X1_261
timestamp 1651764895
transform 1 0 4392 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_382
timestamp 1651764895
transform 1 0 4456 0 -1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_540
timestamp 1651764895
transform 1 0 4488 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_262
timestamp 1651764895
transform 1 0 4552 0 -1 5410
box -4 -6 68 206
use FILL  FILL_26_2_0
timestamp 1651764895
transform 1 0 4616 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_2_1
timestamp 1651764895
transform 1 0 4632 0 -1 5410
box -4 -6 20 206
use FILL  FILL_26_2_2
timestamp 1651764895
transform 1 0 4648 0 -1 5410
box -4 -6 20 206
use NAND3X1  NAND3X1_541
timestamp 1651764895
transform 1 0 4664 0 -1 5410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_84
timestamp 1651764895
transform 1 0 4728 0 -1 5410
box -4 -6 116 206
use AOI21X1  AOI21X1_237
timestamp 1651764895
transform 1 0 4840 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_511
timestamp 1651764895
transform 1 0 4904 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_469
timestamp 1651764895
transform 1 0 4968 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_264
timestamp 1651764895
transform -1 0 5096 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_494
timestamp 1651764895
transform 1 0 5096 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_238
timestamp 1651764895
transform 1 0 5160 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_471
timestamp 1651764895
transform 1 0 5224 0 -1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_470
timestamp 1651764895
transform 1 0 5288 0 -1 5410
box -4 -6 68 206
use INVX1  INVX1_385
timestamp 1651764895
transform 1 0 5352 0 -1 5410
box -4 -6 36 206
use AOI21X1  AOI21X1_266
timestamp 1651764895
transform -1 0 5448 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_499
timestamp 1651764895
transform -1 0 5512 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_503
timestamp 1651764895
transform -1 0 5576 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_489
timestamp 1651764895
transform 1 0 5576 0 -1 5410
box -4 -6 52 206
use NAND3X1  NAND3X1_502
timestamp 1651764895
transform 1 0 5624 0 -1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_240
timestamp 1651764895
transform 1 0 5688 0 -1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_505
timestamp 1651764895
transform -1 0 5816 0 -1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_488
timestamp 1651764895
transform 1 0 5816 0 -1 5410
box -4 -6 52 206
use AOI22X1  AOI22X1_56
timestamp 1651764895
transform 1 0 5864 0 -1 5410
box -4 -6 84 206
use NAND2X1  NAND2X1_544
timestamp 1651764895
transform 1 0 5944 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_14
timestamp 1651764895
transform 1 0 5992 0 -1 5410
box -4 -6 196 206
use NAND2X1  NAND2X1_426
timestamp 1651764895
transform -1 0 6232 0 -1 5410
box -4 -6 52 206
use FILL  FILL_27_1
timestamp 1651764895
transform -1 0 6248 0 -1 5410
box -4 -6 20 206
use FILL  FILL_27_2
timestamp 1651764895
transform -1 0 6264 0 -1 5410
box -4 -6 20 206
use NAND2X1  NAND2X1_522
timestamp 1651764895
transform 1 0 8 0 1 5410
box -4 -6 52 206
use NAND3X1  NAND3X1_517
timestamp 1651764895
transform 1 0 56 0 1 5410
box -4 -6 68 206
use OAI22X1  OAI22X1_12
timestamp 1651764895
transform -1 0 200 0 1 5410
box -4 -6 84 206
use OAI21X1  OAI21X1_494
timestamp 1651764895
transform -1 0 264 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_514
timestamp 1651764895
transform 1 0 264 0 1 5410
box -4 -6 68 206
use OAI22X1  OAI22X1_10
timestamp 1651764895
transform 1 0 328 0 1 5410
box -4 -6 84 206
use NOR2X1  NOR2X1_185
timestamp 1651764895
transform -1 0 456 0 1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_186
timestamp 1651764895
transform 1 0 456 0 1 5410
box -4 -6 52 206
use XNOR2X1  XNOR2X1_67
timestamp 1651764895
transform 1 0 504 0 1 5410
box -4 -6 116 206
use XOR2X1  XOR2X1_45
timestamp 1651764895
transform 1 0 616 0 1 5410
box -4 -6 116 206
use NAND3X1  NAND3X1_519
timestamp 1651764895
transform 1 0 728 0 1 5410
box -4 -6 68 206
use NOR2X1  NOR2X1_184
timestamp 1651764895
transform 1 0 792 0 1 5410
box -4 -6 52 206
use AND2X2  AND2X2_104
timestamp 1651764895
transform -1 0 904 0 1 5410
box -4 -6 68 206
use NOR2X1  NOR2X1_183
timestamp 1651764895
transform -1 0 952 0 1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_182
timestamp 1651764895
transform -1 0 1000 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_435
timestamp 1651764895
transform 1 0 1000 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_456
timestamp 1651764895
transform 1 0 1064 0 1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_181
timestamp 1651764895
transform -1 0 1160 0 1 5410
box -4 -6 52 206
use XOR2X1  XOR2X1_35
timestamp 1651764895
transform -1 0 1272 0 1 5410
box -4 -6 116 206
use OAI21X1  OAI21X1_385
timestamp 1651764895
transform 1 0 1272 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_385
timestamp 1651764895
transform 1 0 1336 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_433
timestamp 1651764895
transform 1 0 1384 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_282
timestamp 1651764895
transform -1 0 1496 0 1 5410
box -4 -6 52 206
use AOI21X1  AOI21X1_197
timestamp 1651764895
transform 1 0 1496 0 1 5410
box -4 -6 68 206
use FILL  FILL_27_0_0
timestamp 1651764895
transform -1 0 1576 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_0_1
timestamp 1651764895
transform -1 0 1592 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_0_2
timestamp 1651764895
transform -1 0 1608 0 1 5410
box -4 -6 20 206
use NOR2X1  NOR2X1_158
timestamp 1651764895
transform -1 0 1656 0 1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_333
timestamp 1651764895
transform 1 0 1656 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_327
timestamp 1651764895
transform 1 0 1704 0 1 5410
box -4 -6 68 206
use XOR2X1  XOR2X1_23
timestamp 1651764895
transform -1 0 1880 0 1 5410
box -4 -6 116 206
use NOR2X1  NOR2X1_139
timestamp 1651764895
transform -1 0 1928 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_382
timestamp 1651764895
transform -1 0 1992 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_309
timestamp 1651764895
transform 1 0 1992 0 1 5410
box -4 -6 36 206
use OR2X2  OR2X2_48
timestamp 1651764895
transform 1 0 2024 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_314
timestamp 1651764895
transform 1 0 2088 0 1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_405
timestamp 1651764895
transform 1 0 2120 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_407
timestamp 1651764895
transform 1 0 2184 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_394
timestamp 1651764895
transform -1 0 2296 0 1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_454
timestamp 1651764895
transform -1 0 2344 0 1 5410
box -4 -6 52 206
use INVX1  INVX1_349
timestamp 1651764895
transform 1 0 2344 0 1 5410
box -4 -6 36 206
use OAI21X1  OAI21X1_497
timestamp 1651764895
transform 1 0 2376 0 1 5410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_48
timestamp 1651764895
transform -1 0 2552 0 1 5410
box -4 -6 116 206
use OR2X2  OR2X2_50
timestamp 1651764895
transform 1 0 2552 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_477
timestamp 1651764895
transform 1 0 2616 0 1 5410
box -4 -6 52 206
use AOI22X1  AOI22X1_53
timestamp 1651764895
transform 1 0 2664 0 1 5410
box -4 -6 84 206
use OAI21X1  OAI21X1_452
timestamp 1651764895
transform 1 0 2744 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_355
timestamp 1651764895
transform -1 0 2840 0 1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_473
timestamp 1651764895
transform 1 0 2840 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_356
timestamp 1651764895
transform -1 0 2936 0 1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_471
timestamp 1651764895
transform 1 0 2936 0 1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_242
timestamp 1651764895
transform 1 0 3000 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_482
timestamp 1651764895
transform 1 0 3064 0 1 5410
box -4 -6 68 206
use FILL  FILL_27_1_0
timestamp 1651764895
transform -1 0 3144 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_1_1
timestamp 1651764895
transform -1 0 3160 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_1_2
timestamp 1651764895
transform -1 0 3176 0 1 5410
box -4 -6 20 206
use AOI21X1  AOI21X1_250
timestamp 1651764895
transform -1 0 3240 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_521
timestamp 1651764895
transform -1 0 3304 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_526
timestamp 1651764895
transform 1 0 3304 0 1 5410
box -4 -6 52 206
use AOI21X1  AOI21X1_251
timestamp 1651764895
transform -1 0 3416 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_523
timestamp 1651764895
transform 1 0 3416 0 1 5410
box -4 -6 68 206
use XOR2X1  XOR2X1_39
timestamp 1651764895
transform 1 0 3480 0 1 5410
box -4 -6 116 206
use NAND2X1  NAND2X1_495
timestamp 1651764895
transform 1 0 3592 0 1 5410
box -4 -6 52 206
use NOR3X1  NOR3X1_47
timestamp 1651764895
transform -1 0 3768 0 1 5410
box -4 -6 132 206
use XOR2X1  XOR2X1_31
timestamp 1651764895
transform -1 0 3880 0 1 5410
box -4 -6 116 206
use NAND2X1  NAND2X1_452
timestamp 1651764895
transform 1 0 3880 0 1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_494
timestamp 1651764895
transform 1 0 3928 0 1 5410
box -4 -6 52 206
use OR2X2  OR2X2_55
timestamp 1651764895
transform 1 0 3976 0 1 5410
box -4 -6 68 206
use AOI22X1  AOI22X1_59
timestamp 1651764895
transform 1 0 4040 0 1 5410
box -4 -6 84 206
use NAND2X1  NAND2X1_541
timestamp 1651764895
transform 1 0 4120 0 1 5410
box -4 -6 52 206
use AND2X2  AND2X2_110
timestamp 1651764895
transform 1 0 4168 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_537
timestamp 1651764895
transform -1 0 4296 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_513
timestamp 1651764895
transform -1 0 4360 0 1 5410
box -4 -6 68 206
use NOR3X1  NOR3X1_51
timestamp 1651764895
transform 1 0 4360 0 1 5410
box -4 -6 132 206
use NAND2X1  NAND2X1_542
timestamp 1651764895
transform 1 0 4488 0 1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_200
timestamp 1651764895
transform -1 0 4584 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_514
timestamp 1651764895
transform 1 0 4584 0 1 5410
box -4 -6 68 206
use FILL  FILL_27_2_0
timestamp 1651764895
transform 1 0 4648 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_2_1
timestamp 1651764895
transform 1 0 4664 0 1 5410
box -4 -6 20 206
use FILL  FILL_27_2_2
timestamp 1651764895
transform 1 0 4680 0 1 5410
box -4 -6 20 206
use NAND3X1  NAND3X1_542
timestamp 1651764895
transform 1 0 4696 0 1 5410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_83
timestamp 1651764895
transform 1 0 4760 0 1 5410
box -4 -6 116 206
use NAND3X1  NAND3X1_543
timestamp 1651764895
transform -1 0 4936 0 1 5410
box -4 -6 68 206
use AOI21X1  AOI21X1_263
timestamp 1651764895
transform 1 0 4936 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_544
timestamp 1651764895
transform -1 0 5064 0 1 5410
box -4 -6 68 206
use AOI22X1  AOI22X1_60
timestamp 1651764895
transform -1 0 5144 0 1 5410
box -4 -6 84 206
use NOR3X1  NOR3X1_52
timestamp 1651764895
transform -1 0 5272 0 1 5410
box -4 -6 132 206
use OAI21X1  OAI21X1_516
timestamp 1651764895
transform 1 0 5272 0 1 5410
box -4 -6 68 206
use INVX1  INVX1_384
timestamp 1651764895
transform 1 0 5336 0 1 5410
box -4 -6 36 206
use AOI21X1  AOI21X1_265
timestamp 1651764895
transform 1 0 5368 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_545
timestamp 1651764895
transform 1 0 5432 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_546
timestamp 1651764895
transform -1 0 5560 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_518
timestamp 1651764895
transform -1 0 5624 0 1 5410
box -4 -6 68 206
use OAI21X1  OAI21X1_515
timestamp 1651764895
transform 1 0 5624 0 1 5410
box -4 -6 68 206
use NAND3X1  NAND3X1_547
timestamp 1651764895
transform 1 0 5688 0 1 5410
box -4 -6 68 206
use NAND2X1  NAND2X1_545
timestamp 1651764895
transform 1 0 5752 0 1 5410
box -4 -6 52 206
use NAND2X1  NAND2X1_543
timestamp 1651764895
transform 1 0 5800 0 1 5410
box -4 -6 52 206
use OAI21X1  OAI21X1_517
timestamp 1651764895
transform -1 0 5912 0 1 5410
box -4 -6 68 206
use NOR2X1  NOR2X1_179
timestamp 1651764895
transform 1 0 5912 0 1 5410
box -4 -6 52 206
use NOR2X1  NOR2X1_178
timestamp 1651764895
transform 1 0 5960 0 1 5410
box -4 -6 52 206
use INVX1  INVX1_386
timestamp 1651764895
transform 1 0 6008 0 1 5410
box -4 -6 36 206
use NAND3X1  NAND3X1_548
timestamp 1651764895
transform 1 0 6040 0 1 5410
box -4 -6 68 206
use BUFX2  BUFX2_31
timestamp 1651764895
transform 1 0 6104 0 1 5410
box -4 -6 52 206
use AOI22X1  AOI22X1_44
timestamp 1651764895
transform 1 0 6152 0 1 5410
box -4 -6 84 206
use FILL  FILL_28_1
timestamp 1651764895
transform 1 0 6232 0 1 5410
box -4 -6 20 206
use FILL  FILL_28_2
timestamp 1651764895
transform 1 0 6248 0 1 5410
box -4 -6 20 206
use NAND3X1  NAND3X1_518
timestamp 1651764895
transform -1 0 72 0 -1 5810
box -4 -6 68 206
use AOI21X1  AOI21X1_246
timestamp 1651764895
transform 1 0 72 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_376
timestamp 1651764895
transform -1 0 168 0 -1 5810
box -4 -6 36 206
use NAND3X1  NAND3X1_516
timestamp 1651764895
transform -1 0 232 0 -1 5810
box -4 -6 68 206
use AOI21X1  AOI21X1_247
timestamp 1651764895
transform 1 0 232 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_495
timestamp 1651764895
transform 1 0 296 0 -1 5810
box -4 -6 68 206
use NAND2X1  NAND2X1_521
timestamp 1651764895
transform -1 0 408 0 -1 5810
box -4 -6 52 206
use NAND3X1  NAND3X1_515
timestamp 1651764895
transform -1 0 472 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_375
timestamp 1651764895
transform -1 0 504 0 -1 5810
box -4 -6 36 206
use INVX1  INVX1_374
timestamp 1651764895
transform 1 0 504 0 -1 5810
box -4 -6 36 206
use OAI21X1  OAI21X1_492
timestamp 1651764895
transform -1 0 600 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_491
timestamp 1651764895
transform -1 0 664 0 -1 5810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_63
timestamp 1651764895
transform 1 0 664 0 -1 5810
box -4 -6 116 206
use NAND2X1  NAND2X1_502
timestamp 1651764895
transform 1 0 776 0 -1 5810
box -4 -6 52 206
use NAND3X1  NAND3X1_462
timestamp 1651764895
transform 1 0 824 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_351
timestamp 1651764895
transform -1 0 920 0 -1 5810
box -4 -6 36 206
use INVX1  INVX1_350
timestamp 1651764895
transform 1 0 920 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_384
timestamp 1651764895
transform -1 0 1000 0 -1 5810
box -4 -6 52 206
use OAI21X1  OAI21X1_434
timestamp 1651764895
transform 1 0 1000 0 -1 5810
box -4 -6 68 206
use NAND2X1  NAND2X1_455
timestamp 1651764895
transform 1 0 1064 0 -1 5810
box -4 -6 52 206
use NAND2X1  NAND2X1_386
timestamp 1651764895
transform 1 0 1112 0 -1 5810
box -4 -6 52 206
use OR2X2  OR2X2_38
timestamp 1651764895
transform -1 0 1224 0 -1 5810
box -4 -6 68 206
use XOR2X1  XOR2X1_27
timestamp 1651764895
transform -1 0 1336 0 -1 5810
box -4 -6 116 206
use NAND2X1  NAND2X1_390
timestamp 1651764895
transform 1 0 1336 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_277
timestamp 1651764895
transform 1 0 1384 0 -1 5810
box -4 -6 36 206
use OAI21X1  OAI21X1_381
timestamp 1651764895
transform -1 0 1480 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_310
timestamp 1651764895
transform -1 0 1512 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_393
timestamp 1651764895
transform 1 0 1512 0 -1 5810
box -4 -6 52 206
use FILL  FILL_28_0_0
timestamp 1651764895
transform -1 0 1576 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_0_1
timestamp 1651764895
transform -1 0 1592 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_0_2
timestamp 1651764895
transform -1 0 1608 0 -1 5810
box -4 -6 20 206
use NAND2X1  NAND2X1_389
timestamp 1651764895
transform -1 0 1656 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_312
timestamp 1651764895
transform -1 0 1688 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_392
timestamp 1651764895
transform 1 0 1688 0 -1 5810
box -4 -6 52 206
use NAND3X1  NAND3X1_403
timestamp 1651764895
transform -1 0 1800 0 -1 5810
box -4 -6 68 206
use AOI21X1  AOI21X1_198
timestamp 1651764895
transform 1 0 1800 0 -1 5810
box -4 -6 68 206
use NAND2X1  NAND2X1_391
timestamp 1651764895
transform 1 0 1864 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_311
timestamp 1651764895
transform -1 0 1944 0 -1 5810
box -4 -6 36 206
use AOI21X1  AOI21X1_199
timestamp 1651764895
transform 1 0 1944 0 -1 5810
box -4 -6 68 206
use NAND3X1  NAND3X1_402
timestamp 1651764895
transform 1 0 2008 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_432
timestamp 1651764895
transform 1 0 2072 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_387
timestamp 1651764895
transform 1 0 2136 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_388
timestamp 1651764895
transform 1 0 2200 0 -1 5810
box -4 -6 68 206
use NAND3X1  NAND3X1_406
timestamp 1651764895
transform 1 0 2264 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_313
timestamp 1651764895
transform -1 0 2360 0 -1 5810
box -4 -6 36 206
use NAND3X1  NAND3X1_404
timestamp 1651764895
transform 1 0 2360 0 -1 5810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_49
timestamp 1651764895
transform 1 0 2424 0 -1 5810
box -4 -6 116 206
use NAND2X1  NAND2X1_460
timestamp 1651764895
transform 1 0 2536 0 -1 5810
box -4 -6 52 206
use NAND3X1  NAND3X1_463
timestamp 1651764895
transform -1 0 2648 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_352
timestamp 1651764895
transform 1 0 2648 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_461
timestamp 1651764895
transform -1 0 2728 0 -1 5810
box -4 -6 52 206
use OAI21X1  OAI21X1_496
timestamp 1651764895
transform 1 0 2728 0 -1 5810
box -4 -6 68 206
use AND2X2  AND2X2_101
timestamp 1651764895
transform 1 0 2792 0 -1 5810
box -4 -6 68 206
use NAND3X1  NAND3X1_467
timestamp 1651764895
transform 1 0 2856 0 -1 5810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_77
timestamp 1651764895
transform 1 0 2920 0 -1 5810
box -4 -6 116 206
use XOR2X1  XOR2X1_50
timestamp 1651764895
transform -1 0 3144 0 -1 5810
box -4 -6 116 206
use FILL  FILL_28_1_0
timestamp 1651764895
transform -1 0 3160 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_1_1
timestamp 1651764895
transform -1 0 3176 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_1_2
timestamp 1651764895
transform -1 0 3192 0 -1 5810
box -4 -6 20 206
use NAND3X1  NAND3X1_520
timestamp 1651764895
transform -1 0 3256 0 -1 5810
box -4 -6 68 206
use NAND2X1  NAND2X1_524
timestamp 1651764895
transform 1 0 3256 0 -1 5810
box -4 -6 52 206
use NAND2X1  NAND2X1_525
timestamp 1651764895
transform 1 0 3304 0 -1 5810
box -4 -6 52 206
use NAND2X1  NAND2X1_523
timestamp 1651764895
transform -1 0 3400 0 -1 5810
box -4 -6 52 206
use NAND3X1  NAND3X1_522
timestamp 1651764895
transform 1 0 3400 0 -1 5810
box -4 -6 68 206
use NOR2X1  NOR2X1_176
timestamp 1651764895
transform -1 0 3512 0 -1 5810
box -4 -6 52 206
use NAND2X1  NAND2X1_485
timestamp 1651764895
transform 1 0 3512 0 -1 5810
box -4 -6 52 206
use OAI21X1  OAI21X1_481
timestamp 1651764895
transform -1 0 3624 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_361
timestamp 1651764895
transform 1 0 3624 0 -1 5810
box -4 -6 36 206
use NOR2X1  NOR2X1_177
timestamp 1651764895
transform -1 0 3704 0 -1 5810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_53
timestamp 1651764895
transform 1 0 3704 0 -1 5810
box -4 -6 116 206
use INVX1  INVX1_360
timestamp 1651764895
transform -1 0 3848 0 -1 5810
box -4 -6 36 206
use OAI21X1  OAI21X1_459
timestamp 1651764895
transform -1 0 3912 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_324
timestamp 1651764895
transform -1 0 3944 0 -1 5810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_45
timestamp 1651764895
transform -1 0 4056 0 -1 5810
box -4 -6 116 206
use NOR2X1  NOR2X1_162
timestamp 1651764895
transform 1 0 4056 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_325
timestamp 1651764895
transform -1 0 4136 0 -1 5810
box -4 -6 36 206
use NOR2X1  NOR2X1_161
timestamp 1651764895
transform 1 0 4136 0 -1 5810
box -4 -6 52 206
use NAND2X1  NAND2X1_415
timestamp 1651764895
transform -1 0 4232 0 -1 5810
box -4 -6 52 206
use XNOR2X1  XNOR2X1_2
timestamp 1651764895
transform 1 0 4232 0 -1 5810
box -4 -6 116 206
use INVX1  INVX1_19
timestamp 1651764895
transform -1 0 4376 0 -1 5810
box -4 -6 36 206
use OAI21X1  OAI21X1_19
timestamp 1651764895
transform 1 0 4376 0 -1 5810
box -4 -6 68 206
use NOR2X1  NOR2X1_20
timestamp 1651764895
transform 1 0 4440 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_20
timestamp 1651764895
transform -1 0 4520 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_14
timestamp 1651764895
transform -1 0 4568 0 -1 5810
box -4 -6 52 206
use NOR2X1  NOR2X1_19
timestamp 1651764895
transform 1 0 4568 0 -1 5810
box -4 -6 52 206
use FILL  FILL_28_2_0
timestamp 1651764895
transform -1 0 4632 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_2_1
timestamp 1651764895
transform -1 0 4648 0 -1 5810
box -4 -6 20 206
use FILL  FILL_28_2_2
timestamp 1651764895
transform -1 0 4664 0 -1 5810
box -4 -6 20 206
use NOR3X1  NOR3X1_48
timestamp 1651764895
transform -1 0 4792 0 -1 5810
box -4 -6 132 206
use OAI21X1  OAI21X1_510
timestamp 1651764895
transform 1 0 4792 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_383
timestamp 1651764895
transform -1 0 4888 0 -1 5810
box -4 -6 36 206
use INVX1  INVX1_381
timestamp 1651764895
transform 1 0 4888 0 -1 5810
box -4 -6 36 206
use INVX1  INVX1_380
timestamp 1651764895
transform 1 0 4920 0 -1 5810
box -4 -6 36 206
use AOI21X1  AOI21X1_259
timestamp 1651764895
transform 1 0 4952 0 -1 5810
box -4 -6 68 206
use NAND3X1  NAND3X1_538
timestamp 1651764895
transform 1 0 5016 0 -1 5810
box -4 -6 68 206
use NAND3X1  NAND3X1_539
timestamp 1651764895
transform -1 0 5144 0 -1 5810
box -4 -6 68 206
use OAI21X1  OAI21X1_509
timestamp 1651764895
transform 1 0 5144 0 -1 5810
box -4 -6 68 206
use INVX1  INVX1_368
timestamp 1651764895
transform -1 0 5240 0 -1 5810
box -4 -6 36 206
use XNOR2X1  XNOR2X1_39
timestamp 1651764895
transform 1 0 5240 0 -1 5810
box -4 -6 116 206
use INVX1  INVX1_292
timestamp 1651764895
transform 1 0 5352 0 -1 5810
box -4 -6 36 206
use OAI21X1  OAI21X1_407
timestamp 1651764895
transform 1 0 5384 0 -1 5810
box -4 -6 68 206
use NOR2X1  NOR2X1_151
timestamp 1651764895
transform 1 0 5448 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_293
timestamp 1651764895
transform -1 0 5528 0 -1 5810
box -4 -6 36 206
use NAND2X1  NAND2X1_354
timestamp 1651764895
transform -1 0 5576 0 -1 5810
box -4 -6 52 206
use NOR2X1  NOR2X1_150
timestamp 1651764895
transform 1 0 5576 0 -1 5810
box -4 -6 52 206
use BUFX2  BUFX2_32
timestamp 1651764895
transform -1 0 5672 0 -1 5810
box -4 -6 52 206
use DFFPOSX1  DFFPOSX1_15
timestamp 1651764895
transform -1 0 5864 0 -1 5810
box -4 -6 196 206
use NAND2X1  NAND2X1_546
timestamp 1651764895
transform -1 0 5912 0 -1 5810
box -4 -6 52 206
use INVX1  INVX1_27
timestamp 1651764895
transform 1 0 5912 0 -1 5810
box -4 -6 36 206
use DFFPOSX1  DFFPOSX1_16
timestamp 1651764895
transform 1 0 5944 0 -1 5810
box -4 -6 196 206
use BUFX2  BUFX2_33
timestamp 1651764895
transform -1 0 6184 0 -1 5810
box -4 -6 52 206
use OAI21X1  OAI21X1_475
timestamp 1651764895
transform -1 0 6248 0 -1 5810
box -4 -6 68 206
use FILL  FILL_29_1
timestamp 1651764895
transform -1 0 6264 0 -1 5810
box -4 -6 20 206
<< labels >>
flabel metal4 s 1560 -40 1608 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 3112 -40 3160 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 5981 5837 5987 5843 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal2 s 493 5837 499 5843 3 FreeSans 24 90 0 0 vertices[0]
port 3 nsew
flabel metal2 s 989 5837 995 5843 3 FreeSans 24 90 0 0 vertices[1]
port 4 nsew
flabel metal2 s 1069 5837 1075 5843 3 FreeSans 24 90 0 0 vertices[2]
port 5 nsew
flabel metal2 s 813 5837 819 5843 3 FreeSans 24 90 0 0 vertices[3]
port 6 nsew
flabel metal3 s -19 1517 -13 1523 7 FreeSans 24 0 0 0 vertices[4]
port 7 nsew
flabel metal3 s -19 2397 -13 2403 7 FreeSans 24 0 0 0 vertices[5]
port 8 nsew
flabel metal3 s -19 2317 -13 2323 7 FreeSans 24 0 0 0 vertices[6]
port 9 nsew
flabel metal3 s -19 2357 -13 2363 7 FreeSans 24 0 0 0 vertices[7]
port 10 nsew
flabel metal3 s -19 2737 -13 2743 7 FreeSans 24 0 0 0 vertices[8]
port 11 nsew
flabel metal3 s -19 4377 -13 4383 7 FreeSans 24 0 0 0 vertices[9]
port 12 nsew
flabel metal3 s -19 3137 -13 3143 7 FreeSans 24 0 0 0 vertices[10]
port 13 nsew
flabel metal3 s -19 3397 -13 3403 7 FreeSans 24 0 0 0 vertices[11]
port 14 nsew
flabel metal3 s -19 3297 -13 3303 7 FreeSans 24 0 0 0 vertices[12]
port 15 nsew
flabel metal3 s -19 3357 -13 3363 7 FreeSans 24 0 0 0 vertices[13]
port 16 nsew
flabel metal3 s -19 3177 -13 3183 7 FreeSans 24 0 0 0 vertices[14]
port 17 nsew
flabel metal3 s -19 2897 -13 2903 7 FreeSans 24 0 0 0 vertices[15]
port 18 nsew
flabel metal3 s -19 2697 -13 2703 7 FreeSans 24 0 0 0 cos_alpha[0]
port 19 nsew
flabel metal3 s -19 2497 -13 2503 7 FreeSans 24 0 0 0 cos_alpha[1]
port 20 nsew
flabel metal3 s -19 1697 -13 1703 7 FreeSans 24 0 0 0 cos_alpha[2]
port 21 nsew
flabel metal3 s -19 3437 -13 3443 7 FreeSans 24 0 0 0 cos_alpha[3]
port 22 nsew
flabel metal3 s -19 3517 -13 3523 7 FreeSans 24 0 0 0 cos_alpha[4]
port 23 nsew
flabel metal3 s -19 4337 -13 4343 7 FreeSans 24 0 0 0 cos_alpha[5]
port 24 nsew
flabel metal3 s -19 4577 -13 4583 7 FreeSans 24 0 0 0 cos_alpha[6]
port 25 nsew
flabel metal3 s -19 3877 -13 3883 7 FreeSans 24 0 0 0 cos_alpha[7]
port 26 nsew
flabel metal3 s -19 4097 -13 4103 7 FreeSans 24 0 0 0 cos_alpha[8]
port 27 nsew
flabel metal2 s 1245 5837 1251 5843 3 FreeSans 24 90 0 0 cos_alpha[9]
port 28 nsew
flabel metal2 s 1469 5837 1475 5843 3 FreeSans 24 90 0 0 cos_alpha[10]
port 29 nsew
flabel metal2 s 1133 5837 1139 5843 3 FreeSans 24 90 0 0 cos_alpha[11]
port 30 nsew
flabel metal2 s 1389 5837 1395 5843 3 FreeSans 24 90 0 0 cos_alpha[12]
port 31 nsew
flabel metal2 s 1501 5837 1507 5843 3 FreeSans 24 90 0 0 cos_alpha[13]
port 32 nsew
flabel metal2 s 925 5837 931 5843 3 FreeSans 24 90 0 0 cos_alpha[14]
port 33 nsew
flabel metal2 s 525 5837 531 5843 3 FreeSans 24 90 0 0 cos_alpha[15]
port 34 nsew
flabel metal3 s -19 2197 -13 2203 7 FreeSans 24 0 0 0 sin_alpha[0]
port 35 nsew
flabel metal2 s 4253 5837 4259 5843 3 FreeSans 24 90 0 0 sin_alpha[1]
port 36 nsew
flabel metal2 s 2077 5837 2083 5843 3 FreeSans 24 90 0 0 sin_alpha[2]
port 37 nsew
flabel metal2 s 877 5837 883 5843 3 FreeSans 24 90 0 0 sin_alpha[3]
port 38 nsew
flabel metal3 s -19 4537 -13 4543 7 FreeSans 24 0 0 0 sin_alpha[4]
port 39 nsew
flabel metal3 s -19 3097 -13 3103 7 FreeSans 24 0 0 0 sin_alpha[5]
port 40 nsew
flabel metal3 s 6285 37 6291 43 3 FreeSans 24 0 0 0 sin_alpha[6]
port 41 nsew
flabel metal3 s -19 3677 -13 3683 7 FreeSans 24 0 0 0 sin_alpha[7]
port 42 nsew
flabel metal3 s 6285 3377 6291 3383 3 FreeSans 24 0 0 0 sin_alpha[8]
port 43 nsew
flabel metal3 s 6285 3417 6291 3423 3 FreeSans 24 0 0 0 sin_alpha[9]
port 44 nsew
flabel metal3 s 6285 4817 6291 4823 3 FreeSans 24 0 0 0 sin_alpha[10]
port 45 nsew
flabel metal3 s -19 5777 -13 5783 7 FreeSans 24 0 0 0 sin_alpha[11]
port 46 nsew
flabel metal3 s 6285 4437 6291 4443 3 FreeSans 24 0 0 0 sin_alpha[12]
port 47 nsew
flabel metal3 s 6285 5237 6291 5243 3 FreeSans 24 0 0 0 sin_alpha[13]
port 48 nsew
flabel metal2 s 1309 -23 1315 -17 7 FreeSans 24 270 0 0 sin_alpha[14]
port 49 nsew
flabel metal3 s -19 5357 -13 5363 7 FreeSans 24 0 0 0 sin_alpha[15]
port 50 nsew
flabel metal3 s 6285 3937 6291 3943 3 FreeSans 24 0 0 0 cos_beta[0]
port 51 nsew
flabel metal3 s 6285 2957 6291 2963 3 FreeSans 24 0 0 0 cos_beta[1]
port 52 nsew
flabel metal3 s -19 5737 -13 5743 7 FreeSans 24 0 0 0 cos_beta[2]
port 53 nsew
flabel metal2 s 1741 5837 1747 5843 3 FreeSans 24 90 0 0 cos_beta[3]
port 54 nsew
flabel metal3 s -19 957 -13 963 7 FreeSans 24 0 0 0 cos_beta[4]
port 55 nsew
flabel metal3 s -19 1817 -13 1823 7 FreeSans 24 0 0 0 cos_beta[5]
port 56 nsew
flabel metal3 s 6285 1137 6291 1143 3 FreeSans 24 0 0 0 cos_beta[6]
port 57 nsew
flabel metal2 s 237 5837 243 5843 3 FreeSans 24 90 0 0 cos_beta[7]
port 58 nsew
flabel metal2 s 2381 5837 2387 5843 3 FreeSans 24 90 0 0 cos_beta[8]
port 59 nsew
flabel metal3 s -19 3777 -13 3783 7 FreeSans 24 0 0 0 cos_beta[9]
port 60 nsew
flabel metal3 s -19 3617 -13 3623 7 FreeSans 24 0 0 0 cos_beta[10]
port 61 nsew
flabel metal3 s 6285 1637 6291 1643 3 FreeSans 24 0 0 0 cos_beta[11]
port 62 nsew
flabel metal3 s -19 1857 -13 1863 7 FreeSans 24 0 0 0 cos_beta[12]
port 63 nsew
flabel metal3 s -19 3557 -13 3563 7 FreeSans 24 0 0 0 cos_beta[13]
port 64 nsew
flabel metal3 s -19 917 -13 923 7 FreeSans 24 0 0 0 cos_beta[14]
port 65 nsew
flabel metal3 s -19 4297 -13 4303 7 FreeSans 24 0 0 0 cos_beta[15]
port 66 nsew
flabel metal2 s 4685 -23 4691 -17 7 FreeSans 24 270 0 0 sin_beta[0]
port 67 nsew
flabel metal2 s 781 5837 787 5843 3 FreeSans 24 90 0 0 sin_beta[1]
port 68 nsew
flabel metal3 s 6285 1777 6291 1783 3 FreeSans 24 0 0 0 sin_beta[2]
port 69 nsew
flabel metal2 s 5005 5837 5011 5843 3 FreeSans 24 90 0 0 sin_beta[3]
port 70 nsew
flabel metal3 s -19 5397 -13 5403 7 FreeSans 24 0 0 0 sin_beta[4]
port 71 nsew
flabel metal3 s -19 37 -13 43 7 FreeSans 24 0 0 0 sin_beta[5]
port 72 nsew
flabel metal3 s -19 3917 -13 3923 7 FreeSans 24 0 0 0 sin_beta[6]
port 73 nsew
flabel metal3 s -19 4797 -13 4803 7 FreeSans 24 0 0 0 sin_beta[7]
port 74 nsew
flabel metal3 s 6285 657 6291 663 3 FreeSans 24 0 0 0 sin_beta[8]
port 75 nsew
flabel metal3 s -19 3057 -13 3063 7 FreeSans 24 0 0 0 sin_beta[9]
port 76 nsew
flabel metal3 s -19 417 -13 423 7 FreeSans 24 0 0 0 sin_beta[10]
port 77 nsew
flabel metal3 s -19 1177 -13 1183 7 FreeSans 24 0 0 0 sin_beta[11]
port 78 nsew
flabel metal3 s 6285 4237 6291 4243 3 FreeSans 24 0 0 0 sin_beta[12]
port 79 nsew
flabel metal2 s 1213 -23 1219 -17 7 FreeSans 24 270 0 0 sin_beta[13]
port 80 nsew
flabel metal2 s 6109 -23 6115 -17 7 FreeSans 24 270 0 0 sin_beta[14]
port 81 nsew
flabel metal3 s 6285 3457 6291 3463 3 FreeSans 24 0 0 0 sin_beta[15]
port 82 nsew
flabel metal2 s 3037 5837 3043 5843 3 FreeSans 24 90 0 0 cos_gamma[0]
port 83 nsew
flabel metal2 s 2781 -23 2787 -17 7 FreeSans 24 270 0 0 cos_gamma[1]
port 84 nsew
flabel metal2 s 2509 -23 2515 -17 7 FreeSans 24 270 0 0 cos_gamma[2]
port 85 nsew
flabel metal2 s 4253 -23 4259 -17 7 FreeSans 24 270 0 0 cos_gamma[3]
port 86 nsew
flabel metal2 s 3437 -23 3443 -17 7 FreeSans 24 270 0 0 cos_gamma[4]
port 87 nsew
flabel metal2 s 4125 -23 4131 -17 7 FreeSans 24 270 0 0 cos_gamma[5]
port 88 nsew
flabel metal2 s 4845 -23 4851 -17 7 FreeSans 24 270 0 0 cos_gamma[6]
port 89 nsew
flabel metal3 s 6285 2997 6291 3003 3 FreeSans 24 0 0 0 cos_gamma[7]
port 90 nsew
flabel metal3 s 6285 2897 6291 2903 3 FreeSans 24 0 0 0 cos_gamma[8]
port 91 nsew
flabel metal3 s 6285 3077 6291 3083 3 FreeSans 24 0 0 0 cos_gamma[9]
port 92 nsew
flabel metal3 s 6285 3037 6291 3043 3 FreeSans 24 0 0 0 cos_gamma[10]
port 93 nsew
flabel metal3 s 6285 3497 6291 3503 3 FreeSans 24 0 0 0 cos_gamma[11]
port 94 nsew
flabel metal3 s 6285 3337 6291 3343 3 FreeSans 24 0 0 0 cos_gamma[12]
port 95 nsew
flabel metal3 s 6285 5297 6291 5303 3 FreeSans 24 0 0 0 cos_gamma[13]
port 96 nsew
flabel metal3 s 6285 317 6291 323 3 FreeSans 24 0 0 0 cos_gamma[14]
port 97 nsew
flabel metal3 s 6285 4097 6291 4103 3 FreeSans 24 0 0 0 cos_gamma[15]
port 98 nsew
flabel metal3 s -19 3977 -13 3983 7 FreeSans 24 0 0 0 sin_gamma[0]
port 99 nsew
flabel metal2 s 5821 5837 5827 5843 3 FreeSans 24 90 0 0 sin_gamma[1]
port 100 nsew
flabel metal2 s 1261 -23 1267 -17 7 FreeSans 24 270 0 0 sin_gamma[2]
port 101 nsew
flabel metal2 s 5869 5837 5875 5843 3 FreeSans 24 90 0 0 sin_gamma[3]
port 102 nsew
flabel metal3 s -19 2777 -13 2783 7 FreeSans 24 0 0 0 sin_gamma[4]
port 103 nsew
flabel metal2 s 4029 5837 4035 5843 3 FreeSans 24 90 0 0 sin_gamma[5]
port 104 nsew
flabel metal2 s 269 5837 275 5843 3 FreeSans 24 90 0 0 sin_gamma[6]
port 105 nsew
flabel metal3 s -19 377 -13 383 7 FreeSans 24 0 0 0 sin_gamma[7]
port 106 nsew
flabel metal2 s 3373 -23 3379 -17 7 FreeSans 24 270 0 0 sin_gamma[8]
port 107 nsew
flabel metal3 s -19 5317 -13 5323 7 FreeSans 24 0 0 0 sin_gamma[9]
port 108 nsew
flabel metal3 s 6285 757 6291 763 3 FreeSans 24 0 0 0 sin_gamma[10]
port 109 nsew
flabel metal2 s 5037 5837 5043 5843 3 FreeSans 24 90 0 0 sin_gamma[11]
port 110 nsew
flabel metal3 s -19 4217 -13 4223 7 FreeSans 24 0 0 0 sin_gamma[12]
port 111 nsew
flabel metal3 s -19 5037 -13 5043 7 FreeSans 24 0 0 0 sin_gamma[13]
port 112 nsew
flabel metal3 s 6285 1897 6291 1903 3 FreeSans 24 0 0 0 sin_gamma[14]
port 113 nsew
flabel metal3 s 6285 2657 6291 2663 3 FreeSans 24 0 0 0 sin_gamma[15]
port 114 nsew
flabel metal2 s 2333 -23 2339 -17 7 FreeSans 24 270 0 0 dx[0]
port 115 nsew
flabel metal2 s 2893 -23 2899 -17 7 FreeSans 24 270 0 0 dx[1]
port 116 nsew
flabel metal2 s 4685 5837 4691 5843 3 FreeSans 24 90 0 0 dx[2]
port 117 nsew
flabel metal2 s 4429 -23 4435 -17 7 FreeSans 24 270 0 0 dx[3]
port 118 nsew
flabel metal2 s 3805 -23 3811 -17 7 FreeSans 24 270 0 0 dx[4]
port 119 nsew
flabel metal2 s 3261 -23 3267 -17 7 FreeSans 24 270 0 0 dx[5]
port 120 nsew
flabel metal2 s 1965 -23 1971 -17 7 FreeSans 24 270 0 0 dx[6]
port 121 nsew
flabel metal2 s 1469 -23 1475 -17 7 FreeSans 24 270 0 0 dx[7]
port 122 nsew
flabel metal2 s 1373 -23 1379 -17 7 FreeSans 24 270 0 0 dx[8]
port 123 nsew
flabel metal2 s 3069 -23 3075 -17 7 FreeSans 24 270 0 0 dx[9]
port 124 nsew
flabel metal2 s 3565 -23 3571 -17 7 FreeSans 24 270 0 0 dx[10]
port 125 nsew
flabel metal3 s 6285 4357 6291 4363 3 FreeSans 24 0 0 0 dx[11]
port 126 nsew
flabel metal2 s 5613 5837 5619 5843 3 FreeSans 24 90 0 0 dx[12]
port 127 nsew
flabel metal2 s 4189 5837 4195 5843 3 FreeSans 24 90 0 0 dx[13]
port 128 nsew
flabel metal2 s 3485 5837 3491 5843 3 FreeSans 24 90 0 0 dx[14]
port 129 nsew
flabel metal3 s 6285 4897 6291 4903 3 FreeSans 24 0 0 0 dx[15]
port 130 nsew
flabel metal2 s 2157 -23 2163 -17 7 FreeSans 24 270 0 0 dy[0]
port 131 nsew
flabel metal2 s 2845 -23 2851 -17 7 FreeSans 24 270 0 0 dy[1]
port 132 nsew
flabel metal2 s 4589 5837 4595 5843 3 FreeSans 24 90 0 0 dy[2]
port 133 nsew
flabel metal2 s 4397 -23 4403 -17 7 FreeSans 24 270 0 0 dy[3]
port 134 nsew
flabel metal2 s 3773 -23 3779 -17 7 FreeSans 24 270 0 0 dy[4]
port 135 nsew
flabel metal2 s 3229 -23 3235 -17 7 FreeSans 24 270 0 0 dy[5]
port 136 nsew
flabel metal2 s 1997 -23 2003 -17 7 FreeSans 24 270 0 0 dy[6]
port 137 nsew
flabel metal2 s 1437 -23 1443 -17 7 FreeSans 24 270 0 0 dy[7]
port 138 nsew
flabel metal2 s 1341 -23 1347 -17 7 FreeSans 24 270 0 0 dy[8]
port 139 nsew
flabel metal2 s 3037 -23 3043 -17 7 FreeSans 24 270 0 0 dy[9]
port 140 nsew
flabel metal2 s 3533 -23 3539 -17 7 FreeSans 24 270 0 0 dy[10]
port 141 nsew
flabel metal3 s 6285 4317 6291 4323 3 FreeSans 24 0 0 0 dy[11]
port 142 nsew
flabel metal2 s 5581 5837 5587 5843 3 FreeSans 24 90 0 0 dy[12]
port 143 nsew
flabel metal2 s 4157 5837 4163 5843 3 FreeSans 24 90 0 0 dy[13]
port 144 nsew
flabel metal2 s 3517 5837 3523 5843 3 FreeSans 24 90 0 0 dy[14]
port 145 nsew
flabel metal2 s 6109 5837 6115 5843 3 FreeSans 24 90 0 0 dy[15]
port 146 nsew
flabel metal2 s 2461 -23 2467 -17 7 FreeSans 24 270 0 0 dz[0]
port 147 nsew
flabel metal2 s 2589 -23 2595 -17 7 FreeSans 24 270 0 0 dz[1]
port 148 nsew
flabel metal2 s 4349 5837 4355 5843 3 FreeSans 24 90 0 0 dz[2]
port 149 nsew
flabel metal2 s 4205 -23 4211 -17 7 FreeSans 24 270 0 0 dz[3]
port 150 nsew
flabel metal2 s 4061 -23 4067 -17 7 FreeSans 24 270 0 0 dz[4]
port 151 nsew
flabel metal2 s 3469 -23 3475 -17 7 FreeSans 24 270 0 0 dz[5]
port 152 nsew
flabel metal2 s 2205 -23 2211 -17 7 FreeSans 24 270 0 0 dz[6]
port 153 nsew
flabel metal2 s 2077 -23 2083 -17 7 FreeSans 24 270 0 0 dz[7]
port 154 nsew
flabel metal2 s 1869 -23 1875 -17 7 FreeSans 24 270 0 0 dz[8]
port 155 nsew
flabel metal2 s 2941 -23 2947 -17 7 FreeSans 24 270 0 0 dz[9]
port 156 nsew
flabel metal2 s 3725 -23 3731 -17 7 FreeSans 24 270 0 0 dz[10]
port 157 nsew
flabel metal3 s 6285 4277 6291 4283 3 FreeSans 24 0 0 0 dz[11]
port 158 nsew
flabel metal2 s 5357 5837 5363 5843 3 FreeSans 24 90 0 0 dz[12]
port 159 nsew
flabel metal2 s 3917 5837 3923 5843 3 FreeSans 24 90 0 0 dz[13]
port 160 nsew
flabel metal2 s 3821 5837 3827 5843 3 FreeSans 24 90 0 0 dz[14]
port 161 nsew
flabel metal3 s 6285 5097 6291 5103 3 FreeSans 24 0 0 0 dz[15]
port 162 nsew
flabel metal2 s 4493 -23 4499 -17 7 FreeSans 24 270 0 0 vertices_out[0]
port 163 nsew
flabel metal2 s 4541 -23 4547 -17 7 FreeSans 24 270 0 0 vertices_out[1]
port 164 nsew
flabel metal3 s 6285 937 6291 943 3 FreeSans 24 0 0 0 vertices_out[2]
port 165 nsew
flabel metal3 s 6285 357 6291 363 3 FreeSans 24 0 0 0 vertices_out[3]
port 166 nsew
flabel metal3 s 6285 897 6291 903 3 FreeSans 24 0 0 0 vertices_out[4]
port 167 nsew
flabel metal2 s 5917 -23 5923 -17 7 FreeSans 24 270 0 0 vertices_out[5]
port 168 nsew
flabel metal2 s 6141 -23 6147 -17 7 FreeSans 24 270 0 0 vertices_out[6]
port 169 nsew
flabel metal2 s 6173 -23 6179 -17 7 FreeSans 24 270 0 0 vertices_out[7]
port 170 nsew
flabel metal3 s 6285 697 6291 703 3 FreeSans 24 0 0 0 vertices_out[8]
port 171 nsew
flabel metal3 s 6285 497 6291 503 3 FreeSans 24 0 0 0 vertices_out[9]
port 172 nsew
flabel metal3 s 6285 1697 6291 1703 3 FreeSans 24 0 0 0 vertices_out[10]
port 173 nsew
flabel metal3 s 6285 2697 6291 2703 3 FreeSans 24 0 0 0 vertices_out[11]
port 174 nsew
flabel metal3 s 6285 3117 6291 3123 3 FreeSans 24 0 0 0 vertices_out[12]
port 175 nsew
flabel metal2 s 6173 5837 6179 5843 3 FreeSans 24 90 0 0 vertices_out[13]
port 176 nsew
flabel metal2 s 5645 5837 5651 5843 3 FreeSans 24 90 0 0 vertices_out[14]
port 177 nsew
flabel metal2 s 6141 5837 6147 5843 3 FreeSans 24 90 0 0 vertices_out[15]
port 178 nsew
<< end >>
